`timescale 1ns / 1ps


module sklanskymod_32_latency_6 (
  input           clk,
  input  [63:0] share0_in,
  input  [63:0] share1_in,
  input  [25:0] rand_bit_share0,
  input  [25:0] rand_bit_share1,
  output [31:0] o_share0,
  output [31:0] o_share1
);

  // Randomness pipeline
  // depth-1 ANDs use rand_bit_share0 directly; deeper ones use these
  wire   [25:0] stage2_share0, stage3_share0, stage4_share0, stage5_share0, stage6_share0;

  reg_26bits rand_stage1 (.clk(clk), .input_share0(rand_bit_share0), .output_share0(stage2_share0));
  reg_26bits rand_stage2 (.clk(clk), .input_share0(stage2_share0), .output_share0(stage3_share0));
  reg_26bits rand_stage3 (.clk(clk), .input_share0(stage3_share0), .output_share0(stage4_share0));
  reg_26bits rand_stage4 (.clk(clk), .input_share0(stage4_share0), .output_share0(stage5_share0));
  reg_26bits rand_stage5 (.clk(clk), .input_share0(stage5_share0), .output_share0(stage6_share0));

  xor_module u_xor_P0_1_d0 (.x_share0(share0_in[1]), .x_share1(share1_in[1]), .y_share0(share0_in[33]), .y_share1(share1_in[33]), .z_share0(d0_P0_1_s0), .z_share1(d0_P0_1_s1));
  xor_module u_xor_P0_10_d0 (.x_share0(share0_in[10]), .x_share1(share1_in[10]), .y_share0(share0_in[42]), .y_share1(share1_in[42]), .z_share0(d0_P0_10_s0), .z_share1(d0_P0_10_s1));
  xor_module u_xor_P0_11_d0 (.x_share0(share0_in[11]), .x_share1(share1_in[11]), .y_share0(share0_in[43]), .y_share1(share1_in[43]), .z_share0(d0_P0_11_s0), .z_share1(d0_P0_11_s1));
  xor_module u_xor_P0_12_d0 (.x_share0(share0_in[12]), .x_share1(share1_in[12]), .y_share0(share0_in[44]), .y_share1(share1_in[44]), .z_share0(d0_P0_12_s0), .z_share1(d0_P0_12_s1));
  xor_module u_xor_P0_13_d0 (.x_share0(share0_in[13]), .x_share1(share1_in[13]), .y_share0(share0_in[45]), .y_share1(share1_in[45]), .z_share0(d0_P0_13_s0), .z_share1(d0_P0_13_s1));
  xor_module u_xor_P0_14_d0 (.x_share0(share0_in[14]), .x_share1(share1_in[14]), .y_share0(share0_in[46]), .y_share1(share1_in[46]), .z_share0(d0_P0_14_s0), .z_share1(d0_P0_14_s1));
  xor_module u_xor_P0_15_d0 (.x_share0(share0_in[15]), .x_share1(share1_in[15]), .y_share0(share0_in[47]), .y_share1(share1_in[47]), .z_share0(d0_P0_15_s0), .z_share1(d0_P0_15_s1));
  xor_module u_xor_P0_16_d0 (.x_share0(share0_in[16]), .x_share1(share1_in[16]), .y_share0(share0_in[48]), .y_share1(share1_in[48]), .z_share0(d0_P0_16_s0), .z_share1(d0_P0_16_s1));
  xor_module u_xor_P0_17_d0 (.x_share0(share0_in[17]), .x_share1(share1_in[17]), .y_share0(share0_in[49]), .y_share1(share1_in[49]), .z_share0(d0_P0_17_s0), .z_share1(d0_P0_17_s1));
  xor_module u_xor_P0_18_d0 (.x_share0(share0_in[18]), .x_share1(share1_in[18]), .y_share0(share0_in[50]), .y_share1(share1_in[50]), .z_share0(d0_P0_18_s0), .z_share1(d0_P0_18_s1));
  xor_module u_xor_P0_19_d0 (.x_share0(share0_in[19]), .x_share1(share1_in[19]), .y_share0(share0_in[51]), .y_share1(share1_in[51]), .z_share0(d0_P0_19_s0), .z_share1(d0_P0_19_s1));
  xor_module u_xor_P0_2_d0 (.x_share0(share0_in[2]), .x_share1(share1_in[2]), .y_share0(share0_in[34]), .y_share1(share1_in[34]), .z_share0(d0_P0_2_s0), .z_share1(d0_P0_2_s1));
  xor_module u_xor_P0_20_d0 (.x_share0(share0_in[20]), .x_share1(share1_in[20]), .y_share0(share0_in[52]), .y_share1(share1_in[52]), .z_share0(d0_P0_20_s0), .z_share1(d0_P0_20_s1));
  xor_module u_xor_P0_21_d0 (.x_share0(share0_in[21]), .x_share1(share1_in[21]), .y_share0(share0_in[53]), .y_share1(share1_in[53]), .z_share0(d0_P0_21_s0), .z_share1(d0_P0_21_s1));
  xor_module u_xor_P0_22_d0 (.x_share0(share0_in[22]), .x_share1(share1_in[22]), .y_share0(share0_in[54]), .y_share1(share1_in[54]), .z_share0(d0_P0_22_s0), .z_share1(d0_P0_22_s1));
  xor_module u_xor_P0_23_d0 (.x_share0(share0_in[23]), .x_share1(share1_in[23]), .y_share0(share0_in[55]), .y_share1(share1_in[55]), .z_share0(d0_P0_23_s0), .z_share1(d0_P0_23_s1));
  xor_module u_xor_P0_24_d0 (.x_share0(share0_in[24]), .x_share1(share1_in[24]), .y_share0(share0_in[56]), .y_share1(share1_in[56]), .z_share0(d0_P0_24_s0), .z_share1(d0_P0_24_s1));
  xor_module u_xor_P0_25_d0 (.x_share0(share0_in[25]), .x_share1(share1_in[25]), .y_share0(share0_in[57]), .y_share1(share1_in[57]), .z_share0(d0_P0_25_s0), .z_share1(d0_P0_25_s1));
  xor_module u_xor_P0_26_d0 (.x_share0(share0_in[26]), .x_share1(share1_in[26]), .y_share0(share0_in[58]), .y_share1(share1_in[58]), .z_share0(d0_P0_26_s0), .z_share1(d0_P0_26_s1));
  xor_module u_xor_P0_27_d0 (.x_share0(share0_in[27]), .x_share1(share1_in[27]), .y_share0(share0_in[59]), .y_share1(share1_in[59]), .z_share0(d0_P0_27_s0), .z_share1(d0_P0_27_s1));
  xor_module u_xor_P0_28_d0 (.x_share0(share0_in[28]), .x_share1(share1_in[28]), .y_share0(share0_in[60]), .y_share1(share1_in[60]), .z_share0(d0_P0_28_s0), .z_share1(d0_P0_28_s1));
  xor_module u_xor_P0_29_d0 (.x_share0(share0_in[29]), .x_share1(share1_in[29]), .y_share0(share0_in[61]), .y_share1(share1_in[61]), .z_share0(d0_P0_29_s0), .z_share1(d0_P0_29_s1));
  xor_module u_xor_P0_3_d0 (.x_share0(share0_in[3]), .x_share1(share1_in[3]), .y_share0(share0_in[35]), .y_share1(share1_in[35]), .z_share0(d0_P0_3_s0), .z_share1(d0_P0_3_s1));
  xor_module u_xor_P0_30_d0 (.x_share0(share0_in[30]), .x_share1(share1_in[30]), .y_share0(share0_in[62]), .y_share1(share1_in[62]), .z_share0(d0_P0_30_s0), .z_share1(d0_P0_30_s1));
  xor_module u_xor_P0_31_d0 (.x_share0(share0_in[31]), .x_share1(share1_in[31]), .y_share0(share0_in[63]), .y_share1(share1_in[63]), .z_share0(d0_P0_31_s0), .z_share1(d0_P0_31_s1));
  xor_module u_xor_P0_4_d0 (.x_share0(share0_in[4]), .x_share1(share1_in[4]), .y_share0(share0_in[36]), .y_share1(share1_in[36]), .z_share0(d0_P0_4_s0), .z_share1(d0_P0_4_s1));
  xor_module u_xor_P0_5_d0 (.x_share0(share0_in[5]), .x_share1(share1_in[5]), .y_share0(share0_in[37]), .y_share1(share1_in[37]), .z_share0(d0_P0_5_s0), .z_share1(d0_P0_5_s1));
  xor_module u_xor_P0_6_d0 (.x_share0(share0_in[6]), .x_share1(share1_in[6]), .y_share0(share0_in[38]), .y_share1(share1_in[38]), .z_share0(d0_P0_6_s0), .z_share1(d0_P0_6_s1));
  xor_module u_xor_P0_7_d0 (.x_share0(share0_in[7]), .x_share1(share1_in[7]), .y_share0(share0_in[39]), .y_share1(share1_in[39]), .z_share0(d0_P0_7_s0), .z_share1(d0_P0_7_s1));
  xor_module u_xor_P0_8_d0 (.x_share0(share0_in[8]), .x_share1(share1_in[8]), .y_share0(share0_in[40]), .y_share1(share1_in[40]), .z_share0(d0_P0_8_s0), .z_share1(d0_P0_8_s1));
  xor_module u_xor_P0_9_d0 (.x_share0(share0_in[9]), .x_share1(share1_in[9]), .y_share0(share0_in[41]), .y_share1(share1_in[41]), .z_share0(d0_P0_9_s0), .z_share1(d0_P0_9_s1));
  xor_module u_xor_o0_d0 (.x_share0(share0_in[0]), .x_share1(share1_in[0]), .y_share0(share0_in[32]), .y_share1(share1_in[32]), .z_share0(d0_o0_s0), .z_share1(d0_o0_s1));
  reg_module u_reg_P0_1_d1 (.clk(clk), .input_share0(d0_P0_1_s0), .input_share1(d0_P0_1_s1), .output_share0(d1_P0_1_s0), .output_share1(d1_P0_1_s1));
  reg_module u_reg_P0_10_d1 (.clk(clk), .input_share0(d0_P0_10_s0), .input_share1(d0_P0_10_s1), .output_share0(d1_P0_10_s0), .output_share1(d1_P0_10_s1));
  reg_module u_reg_P0_11_d1 (.clk(clk), .input_share0(d0_P0_11_s0), .input_share1(d0_P0_11_s1), .output_share0(d1_P0_11_s0), .output_share1(d1_P0_11_s1));
  reg_module u_reg_P0_12_d1 (.clk(clk), .input_share0(d0_P0_12_s0), .input_share1(d0_P0_12_s1), .output_share0(d1_P0_12_s0), .output_share1(d1_P0_12_s1));
  reg_module u_reg_P0_13_d1 (.clk(clk), .input_share0(d0_P0_13_s0), .input_share1(d0_P0_13_s1), .output_share0(d1_P0_13_s0), .output_share1(d1_P0_13_s1));
  reg_module u_reg_P0_14_d1 (.clk(clk), .input_share0(d0_P0_14_s0), .input_share1(d0_P0_14_s1), .output_share0(d1_P0_14_s0), .output_share1(d1_P0_14_s1));
  reg_module u_reg_P0_15_d1 (.clk(clk), .input_share0(d0_P0_15_s0), .input_share1(d0_P0_15_s1), .output_share0(d1_P0_15_s0), .output_share1(d1_P0_15_s1));
  reg_module u_reg_P0_16_d1 (.clk(clk), .input_share0(d0_P0_16_s0), .input_share1(d0_P0_16_s1), .output_share0(d1_P0_16_s0), .output_share1(d1_P0_16_s1));
  reg_module u_reg_P0_17_d1 (.clk(clk), .input_share0(d0_P0_17_s0), .input_share1(d0_P0_17_s1), .output_share0(d1_P0_17_s0), .output_share1(d1_P0_17_s1));
  reg_module u_reg_P0_18_d1 (.clk(clk), .input_share0(d0_P0_18_s0), .input_share1(d0_P0_18_s1), .output_share0(d1_P0_18_s0), .output_share1(d1_P0_18_s1));
  reg_module u_reg_P0_19_d1 (.clk(clk), .input_share0(d0_P0_19_s0), .input_share1(d0_P0_19_s1), .output_share0(d1_P0_19_s0), .output_share1(d1_P0_19_s1));
  reg_module u_reg_P0_2_d1 (.clk(clk), .input_share0(d0_P0_2_s0), .input_share1(d0_P0_2_s1), .output_share0(d1_P0_2_s0), .output_share1(d1_P0_2_s1));
  reg_module u_reg_P0_20_d1 (.clk(clk), .input_share0(d0_P0_20_s0), .input_share1(d0_P0_20_s1), .output_share0(d1_P0_20_s0), .output_share1(d1_P0_20_s1));
  reg_module u_reg_P0_21_d1 (.clk(clk), .input_share0(d0_P0_21_s0), .input_share1(d0_P0_21_s1), .output_share0(d1_P0_21_s0), .output_share1(d1_P0_21_s1));
  reg_module u_reg_P0_22_d1 (.clk(clk), .input_share0(d0_P0_22_s0), .input_share1(d0_P0_22_s1), .output_share0(d1_P0_22_s0), .output_share1(d1_P0_22_s1));
  reg_module u_reg_P0_23_d1 (.clk(clk), .input_share0(d0_P0_23_s0), .input_share1(d0_P0_23_s1), .output_share0(d1_P0_23_s0), .output_share1(d1_P0_23_s1));
  reg_module u_reg_P0_24_d1 (.clk(clk), .input_share0(d0_P0_24_s0), .input_share1(d0_P0_24_s1), .output_share0(d1_P0_24_s0), .output_share1(d1_P0_24_s1));
  reg_module u_reg_P0_25_d1 (.clk(clk), .input_share0(d0_P0_25_s0), .input_share1(d0_P0_25_s1), .output_share0(d1_P0_25_s0), .output_share1(d1_P0_25_s1));
  reg_module u_reg_P0_26_d1 (.clk(clk), .input_share0(d0_P0_26_s0), .input_share1(d0_P0_26_s1), .output_share0(d1_P0_26_s0), .output_share1(d1_P0_26_s1));
  reg_module u_reg_P0_27_d1 (.clk(clk), .input_share0(d0_P0_27_s0), .input_share1(d0_P0_27_s1), .output_share0(d1_P0_27_s0), .output_share1(d1_P0_27_s1));
  reg_module u_reg_P0_28_d1 (.clk(clk), .input_share0(d0_P0_28_s0), .input_share1(d0_P0_28_s1), .output_share0(d1_P0_28_s0), .output_share1(d1_P0_28_s1));
  reg_module u_reg_P0_29_d1 (.clk(clk), .input_share0(d0_P0_29_s0), .input_share1(d0_P0_29_s1), .output_share0(d1_P0_29_s0), .output_share1(d1_P0_29_s1));
  reg_module u_reg_P0_3_d1 (.clk(clk), .input_share0(d0_P0_3_s0), .input_share1(d0_P0_3_s1), .output_share0(d1_P0_3_s0), .output_share1(d1_P0_3_s1));
  reg_module u_reg_P0_30_d1 (.clk(clk), .input_share0(d0_P0_30_s0), .input_share1(d0_P0_30_s1), .output_share0(d1_P0_30_s0), .output_share1(d1_P0_30_s1));
  reg_module u_reg_P0_31_d1 (.clk(clk), .input_share0(d0_P0_31_s0), .input_share1(d0_P0_31_s1), .output_share0(d1_P0_31_s0), .output_share1(d1_P0_31_s1));
  reg_module u_reg_P0_4_d1 (.clk(clk), .input_share0(d0_P0_4_s0), .input_share1(d0_P0_4_s1), .output_share0(d1_P0_4_s0), .output_share1(d1_P0_4_s1));
  reg_module u_reg_P0_5_d1 (.clk(clk), .input_share0(d0_P0_5_s0), .input_share1(d0_P0_5_s1), .output_share0(d1_P0_5_s0), .output_share1(d1_P0_5_s1));
  reg_module u_reg_P0_6_d1 (.clk(clk), .input_share0(d0_P0_6_s0), .input_share1(d0_P0_6_s1), .output_share0(d1_P0_6_s0), .output_share1(d1_P0_6_s1));
  reg_module u_reg_P0_7_d1 (.clk(clk), .input_share0(d0_P0_7_s0), .input_share1(d0_P0_7_s1), .output_share0(d1_P0_7_s0), .output_share1(d1_P0_7_s1));
  reg_module u_reg_P0_8_d1 (.clk(clk), .input_share0(d0_P0_8_s0), .input_share1(d0_P0_8_s1), .output_share0(d1_P0_8_s0), .output_share1(d1_P0_8_s1));
  reg_module u_reg_P0_9_d1 (.clk(clk), .input_share0(d0_P0_9_s0), .input_share1(d0_P0_9_s1), .output_share0(d1_P0_9_s0), .output_share1(d1_P0_9_s1));
  and_module u_and_G0_0_d1 (.clk(clk), .x_share0(share0_in[0]), .x_share1(share1_in[0]), .y_share0(share0_in[32]), .y_share1(share1_in[32]), .rand(r_G0_0), .z_share0(d1_G0_0_s0), .z_share1(d1_G0_0_s1));
  assign r_G0_0 = rand_bit_share0[2];
  and_module u_and_G0_1_d1 (.clk(clk), .x_share0(share0_in[1]), .x_share1(share1_in[1]), .y_share0(share0_in[33]), .y_share1(share1_in[33]), .rand(r_G0_1), .z_share0(d1_G0_1_s0), .z_share1(d1_G0_1_s1));
  assign r_G0_1 = rand_bit_share0[0];
  and_module u_and_G0_10_d1 (.clk(clk), .x_share0(share0_in[10]), .x_share1(share1_in[10]), .y_share0(share0_in[42]), .y_share1(share1_in[42]), .rand(r_G0_10), .z_share0(d1_G0_10_s0), .z_share1(d1_G0_10_s1));
  assign r_G0_10 = rand_bit_share0[1];
  and_module u_and_G0_11_d1 (.clk(clk), .x_share0(share0_in[11]), .x_share1(share1_in[11]), .y_share0(share0_in[43]), .y_share1(share1_in[43]), .rand(r_G0_11), .z_share0(d1_G0_11_s0), .z_share1(d1_G0_11_s1));
  assign r_G0_11 = rand_bit_share0[2];
  and_module u_and_G0_12_d1 (.clk(clk), .x_share0(share0_in[12]), .x_share1(share1_in[12]), .y_share0(share0_in[44]), .y_share1(share1_in[44]), .rand(r_G0_12), .z_share0(d1_G0_12_s0), .z_share1(d1_G0_12_s1));
  assign r_G0_12 = rand_bit_share0[3];
  and_module u_and_G0_13_d1 (.clk(clk), .x_share0(share0_in[13]), .x_share1(share1_in[13]), .y_share0(share0_in[45]), .y_share1(share1_in[45]), .rand(r_G0_13), .z_share0(d1_G0_13_s0), .z_share1(d1_G0_13_s1));
  assign r_G0_13 = rand_bit_share0[1];
  and_module u_and_G0_14_d1 (.clk(clk), .x_share0(share0_in[14]), .x_share1(share1_in[14]), .y_share0(share0_in[46]), .y_share1(share1_in[46]), .rand(r_G0_14), .z_share0(d1_G0_14_s0), .z_share1(d1_G0_14_s1));
  assign r_G0_14 = rand_bit_share0[0];
  and_module u_and_G0_15_d1 (.clk(clk), .x_share0(share0_in[15]), .x_share1(share1_in[15]), .y_share0(share0_in[47]), .y_share1(share1_in[47]), .rand(r_G0_15), .z_share0(d1_G0_15_s0), .z_share1(d1_G0_15_s1));
  assign r_G0_15 = rand_bit_share0[3];
  and_module u_and_G0_16_d1 (.clk(clk), .x_share0(share0_in[16]), .x_share1(share1_in[16]), .y_share0(share0_in[48]), .y_share1(share1_in[48]), .rand(r_G0_16), .z_share0(d1_G0_16_s0), .z_share1(d1_G0_16_s1));
  assign r_G0_16 = rand_bit_share0[10];
  and_module u_and_G0_17_d1 (.clk(clk), .x_share0(share0_in[17]), .x_share1(share1_in[17]), .y_share0(share0_in[49]), .y_share1(share1_in[49]), .rand(r_G0_17), .z_share0(d1_G0_17_s0), .z_share1(d1_G0_17_s1));
  assign r_G0_17 = rand_bit_share0[8];
  and_module u_and_G0_18_d1 (.clk(clk), .x_share0(share0_in[18]), .x_share1(share1_in[18]), .y_share0(share0_in[50]), .y_share1(share1_in[50]), .rand(r_G0_18), .z_share0(d1_G0_18_s0), .z_share1(d1_G0_18_s1));
  assign r_G0_18 = rand_bit_share0[10];
  and_module u_and_G0_19_d1 (.clk(clk), .x_share0(share0_in[19]), .x_share1(share1_in[19]), .y_share0(share0_in[51]), .y_share1(share1_in[51]), .rand(r_G0_19), .z_share0(d1_G0_19_s0), .z_share1(d1_G0_19_s1));
  assign r_G0_19 = rand_bit_share0[12];
  and_module u_and_G0_2_d1 (.clk(clk), .x_share0(share0_in[2]), .x_share1(share1_in[2]), .y_share0(share0_in[34]), .y_share1(share1_in[34]), .rand(r_G0_2), .z_share0(d1_G0_2_s0), .z_share1(d1_G0_2_s1));
  assign r_G0_2 = rand_bit_share0[2];
  and_module u_and_G0_20_d1 (.clk(clk), .x_share0(share0_in[20]), .x_share1(share1_in[20]), .y_share0(share0_in[52]), .y_share1(share1_in[52]), .rand(r_G0_20), .z_share0(d1_G0_20_s0), .z_share1(d1_G0_20_s1));
  assign r_G0_20 = rand_bit_share0[8];
  and_module u_and_G0_21_d1 (.clk(clk), .x_share0(share0_in[21]), .x_share1(share1_in[21]), .y_share0(share0_in[53]), .y_share1(share1_in[53]), .rand(r_G0_21), .z_share0(d1_G0_21_s0), .z_share1(d1_G0_21_s1));
  assign r_G0_21 = rand_bit_share0[11];
  and_module u_and_G0_22_d1 (.clk(clk), .x_share0(share0_in[22]), .x_share1(share1_in[22]), .y_share0(share0_in[54]), .y_share1(share1_in[54]), .rand(r_G0_22), .z_share0(d1_G0_22_s0), .z_share1(d1_G0_22_s1));
  assign r_G0_22 = rand_bit_share0[10];
  and_module u_and_G0_23_d1 (.clk(clk), .x_share0(share0_in[23]), .x_share1(share1_in[23]), .y_share0(share0_in[55]), .y_share1(share1_in[55]), .rand(r_G0_23), .z_share0(d1_G0_23_s0), .z_share1(d1_G0_23_s1));
  assign r_G0_23 = rand_bit_share0[8];
  and_module u_and_G0_24_d1 (.clk(clk), .x_share0(share0_in[24]), .x_share1(share1_in[24]), .y_share0(share0_in[56]), .y_share1(share1_in[56]), .rand(r_G0_24), .z_share0(d1_G0_24_s0), .z_share1(d1_G0_24_s1));
  assign r_G0_24 = rand_bit_share0[13];
  and_module u_and_G0_25_d1 (.clk(clk), .x_share0(share0_in[25]), .x_share1(share1_in[25]), .y_share0(share0_in[57]), .y_share1(share1_in[57]), .rand(r_G0_25), .z_share0(d1_G0_25_s0), .z_share1(d1_G0_25_s1));
  assign r_G0_25 = rand_bit_share0[18];
  and_module u_and_G0_26_d1 (.clk(clk), .x_share0(share0_in[26]), .x_share1(share1_in[26]), .y_share0(share0_in[58]), .y_share1(share1_in[58]), .rand(r_G0_26), .z_share0(d1_G0_26_s0), .z_share1(d1_G0_26_s1));
  assign r_G0_26 = rand_bit_share0[16];
  and_module u_and_G0_27_d1 (.clk(clk), .x_share0(share0_in[27]), .x_share1(share1_in[27]), .y_share0(share0_in[59]), .y_share1(share1_in[59]), .rand(r_G0_27), .z_share0(d1_G0_27_s0), .z_share1(d1_G0_27_s1));
  assign r_G0_27 = rand_bit_share0[12];
  and_module u_and_G0_28_d1 (.clk(clk), .x_share0(share0_in[28]), .x_share1(share1_in[28]), .y_share0(share0_in[60]), .y_share1(share1_in[60]), .rand(r_G0_28), .z_share0(d1_G0_28_s0), .z_share1(d1_G0_28_s1));
  assign r_G0_28 = rand_bit_share0[21];
  and_module u_and_G0_29_d1 (.clk(clk), .x_share0(share0_in[29]), .x_share1(share1_in[29]), .y_share0(share0_in[61]), .y_share1(share1_in[61]), .rand(r_G0_29), .z_share0(d1_G0_29_s0), .z_share1(d1_G0_29_s1));
  assign r_G0_29 = rand_bit_share0[22];
  and_module u_and_G0_3_d1 (.clk(clk), .x_share0(share0_in[3]), .x_share1(share1_in[3]), .y_share0(share0_in[35]), .y_share1(share1_in[35]), .rand(r_G0_3), .z_share0(d1_G0_3_s0), .z_share1(d1_G0_3_s1));
  assign r_G0_3 = rand_bit_share0[5];
  and_module u_and_G0_30_d1 (.clk(clk), .x_share0(share0_in[30]), .x_share1(share1_in[30]), .y_share0(share0_in[62]), .y_share1(share1_in[62]), .rand(r_G0_30), .z_share0(d1_G0_30_s0), .z_share1(d1_G0_30_s1));
  assign r_G0_30 = rand_bit_share0[24];
  and_module u_and_G0_31_d1 (.clk(clk), .x_share0(share0_in[31]), .x_share1(share1_in[31]), .y_share0(share0_in[63]), .y_share1(share1_in[63]), .rand(r_G0_31), .z_share0(d1_G0_31_s0), .z_share1(d1_G0_31_s1));
  assign r_G0_31 = rand_bit_share0[18];
  and_module u_and_G0_4_d1 (.clk(clk), .x_share0(share0_in[4]), .x_share1(share1_in[4]), .y_share0(share0_in[36]), .y_share1(share1_in[36]), .rand(r_G0_4), .z_share0(d1_G0_4_s0), .z_share1(d1_G0_4_s1));
  assign r_G0_4 = rand_bit_share0[2];
  and_module u_and_G0_5_d1 (.clk(clk), .x_share0(share0_in[5]), .x_share1(share1_in[5]), .y_share0(share0_in[37]), .y_share1(share1_in[37]), .rand(r_G0_5), .z_share0(d1_G0_5_s0), .z_share1(d1_G0_5_s1));
  assign r_G0_5 = rand_bit_share0[0];
  and_module u_and_G0_6_d1 (.clk(clk), .x_share0(share0_in[6]), .x_share1(share1_in[6]), .y_share0(share0_in[38]), .y_share1(share1_in[38]), .rand(r_G0_6), .z_share0(d1_G0_6_s0), .z_share1(d1_G0_6_s1));
  assign r_G0_6 = rand_bit_share0[2];
  and_module u_and_G0_7_d1 (.clk(clk), .x_share0(share0_in[7]), .x_share1(share1_in[7]), .y_share0(share0_in[39]), .y_share1(share1_in[39]), .rand(r_G0_7), .z_share0(d1_G0_7_s0), .z_share1(d1_G0_7_s1));
  assign r_G0_7 = rand_bit_share0[9];
  and_module u_and_G0_8_d1 (.clk(clk), .x_share0(share0_in[8]), .x_share1(share1_in[8]), .y_share0(share0_in[40]), .y_share1(share1_in[40]), .rand(r_G0_8), .z_share0(d1_G0_8_s0), .z_share1(d1_G0_8_s1));
  assign r_G0_8 = rand_bit_share0[0];
  and_module u_and_G0_9_d1 (.clk(clk), .x_share0(share0_in[9]), .x_share1(share1_in[9]), .y_share0(share0_in[41]), .y_share1(share1_in[41]), .rand(r_G0_9), .z_share0(d1_G0_9_s0), .z_share1(d1_G0_9_s1));
  assign r_G0_9 = rand_bit_share0[4];
  and_module u_and_P1_11_d1 (.clk(clk), .x_share0(d0_P0_11_s0), .x_share1(d0_P0_11_s1), .y_share0(d0_P0_10_s0), .y_share1(d0_P0_10_s1), .rand(r_P1_11), .z_share0(d1_P1_11_s0), .z_share1(d1_P1_11_s1));
  assign r_P1_11 = rand_bit_share0[7];
  and_module u_and_P1_13_d1 (.clk(clk), .x_share0(d0_P0_13_s0), .x_share1(d0_P0_13_s1), .y_share0(d0_P0_12_s0), .y_share1(d0_P0_12_s1), .rand(r_P1_13), .z_share0(d1_P1_13_s0), .z_share1(d1_P1_13_s1));
  assign r_P1_13 = rand_bit_share0[3];
  and_module u_and_P1_15_d1 (.clk(clk), .x_share0(d0_P0_15_s0), .x_share1(d0_P0_15_s1), .y_share0(d0_P0_14_s0), .y_share1(d0_P0_14_s1), .rand(r_P1_15), .z_share0(d1_P1_15_s0), .z_share1(d1_P1_15_s1));
  assign r_P1_15 = rand_bit_share0[0];
  and_module u_and_P1_17_d1 (.clk(clk), .x_share0(d0_P0_17_s0), .x_share1(d0_P0_17_s1), .y_share0(d0_P0_16_s0), .y_share1(d0_P0_16_s1), .rand(r_P1_17), .z_share0(d1_P1_17_s0), .z_share1(d1_P1_17_s1));
  assign r_P1_17 = rand_bit_share0[19];
  and_module u_and_P1_19_d1 (.clk(clk), .x_share0(d0_P0_19_s0), .x_share1(d0_P0_19_s1), .y_share0(d0_P0_18_s0), .y_share1(d0_P0_18_s1), .rand(r_P1_19), .z_share0(d1_P1_19_s0), .z_share1(d1_P1_19_s1));
  assign r_P1_19 = rand_bit_share0[16];
  and_module u_and_P1_21_d1 (.clk(clk), .x_share0(d0_P0_21_s0), .x_share1(d0_P0_21_s1), .y_share0(d0_P0_20_s0), .y_share1(d0_P0_20_s1), .rand(r_P1_21), .z_share0(d1_P1_21_s0), .z_share1(d1_P1_21_s1));
  assign r_P1_21 = rand_bit_share0[17];
  and_module u_and_P1_23_d1 (.clk(clk), .x_share0(d0_P0_23_s0), .x_share1(d0_P0_23_s1), .y_share0(d0_P0_22_s0), .y_share1(d0_P0_22_s1), .rand(r_P1_23), .z_share0(d1_P1_23_s0), .z_share1(d1_P1_23_s1));
  assign r_P1_23 = rand_bit_share0[14];
  and_module u_and_P1_25_d1 (.clk(clk), .x_share0(d0_P0_25_s0), .x_share1(d0_P0_25_s1), .y_share0(d0_P0_24_s0), .y_share1(d0_P0_24_s1), .rand(r_P1_25), .z_share0(d1_P1_25_s0), .z_share1(d1_P1_25_s1));
  assign r_P1_25 = rand_bit_share0[24];
  and_module u_and_P1_27_d1 (.clk(clk), .x_share0(d0_P0_27_s0), .x_share1(d0_P0_27_s1), .y_share0(d0_P0_26_s0), .y_share1(d0_P0_26_s1), .rand(r_P1_27), .z_share0(d1_P1_27_s0), .z_share1(d1_P1_27_s1));
  assign r_P1_27 = rand_bit_share0[17];
  and_module u_and_P1_29_d1 (.clk(clk), .x_share0(d0_P0_29_s0), .x_share1(d0_P0_29_s1), .y_share0(d0_P0_28_s0), .y_share1(d0_P0_28_s1), .rand(r_P1_29), .z_share0(d1_P1_29_s0), .z_share1(d1_P1_29_s1));
  assign r_P1_29 = rand_bit_share0[20];
  and_module u_and_P1_3_d1 (.clk(clk), .x_share0(d0_P0_3_s0), .x_share1(d0_P0_3_s1), .y_share0(d0_P0_2_s0), .y_share1(d0_P0_2_s1), .rand(r_P1_3), .z_share0(d1_P1_3_s0), .z_share1(d1_P1_3_s1));
  assign r_P1_3 = rand_bit_share0[14];
  and_module u_and_P1_31_d1 (.clk(clk), .x_share0(d0_P0_31_s0), .x_share1(d0_P0_31_s1), .y_share0(d0_P0_30_s0), .y_share1(d0_P0_30_s1), .rand(r_P1_31), .z_share0(d1_P1_31_s0), .z_share1(d1_P1_31_s1));
  assign r_P1_31 = rand_bit_share0[19];
  and_module u_and_P1_5_d1 (.clk(clk), .x_share0(d0_P0_5_s0), .x_share1(d0_P0_5_s1), .y_share0(d0_P0_4_s0), .y_share1(d0_P0_4_s1), .rand(r_P1_5), .z_share0(d1_P1_5_s0), .z_share1(d1_P1_5_s1));
  assign r_P1_5 = rand_bit_share0[2];
  and_module u_and_P1_7_d1 (.clk(clk), .x_share0(d0_P0_7_s0), .x_share1(d0_P0_7_s1), .y_share0(d0_P0_6_s0), .y_share1(d0_P0_6_s1), .rand(r_P1_7), .z_share0(d1_P1_7_s0), .z_share1(d1_P1_7_s1));
  assign r_P1_7 = rand_bit_share0[8];
  and_module u_and_P1_9_d1 (.clk(clk), .x_share0(d0_P0_9_s0), .x_share1(d0_P0_9_s1), .y_share0(d0_P0_8_s0), .y_share1(d0_P0_8_s1), .rand(r_P1_9), .z_share0(d1_P1_9_s0), .z_share1(d1_P1_9_s1));
  assign r_P1_9 = rand_bit_share0[6];
  xor_module u_xor_o1_d1 (.x_share0(d1_P0_1_s0), .x_share1(d1_P0_1_s1), .y_share0(d1_G0_0_s0), .y_share1(d1_G0_0_s1), .z_share0(d1_o1_s0), .z_share1(d1_o1_s1));
  reg_module u_reg_G0_1_d2 (.clk(clk), .input_share0(d1_G0_1_s0), .input_share1(d1_G0_1_s1), .output_share0(d2_G0_1_s0), .output_share1(d2_G0_1_s1));
  reg_module u_reg_G0_10_d2 (.clk(clk), .input_share0(d1_G0_10_s0), .input_share1(d1_G0_10_s1), .output_share0(d2_G0_10_s0), .output_share1(d2_G0_10_s1));
  reg_module u_reg_G0_11_d2 (.clk(clk), .input_share0(d1_G0_11_s0), .input_share1(d1_G0_11_s1), .output_share0(d2_G0_11_s0), .output_share1(d2_G0_11_s1));
  reg_module u_reg_G0_12_d2 (.clk(clk), .input_share0(d1_G0_12_s0), .input_share1(d1_G0_12_s1), .output_share0(d2_G0_12_s0), .output_share1(d2_G0_12_s1));
  reg_module u_reg_G0_13_d2 (.clk(clk), .input_share0(d1_G0_13_s0), .input_share1(d1_G0_13_s1), .output_share0(d2_G0_13_s0), .output_share1(d2_G0_13_s1));
  reg_module u_reg_G0_14_d2 (.clk(clk), .input_share0(d1_G0_14_s0), .input_share1(d1_G0_14_s1), .output_share0(d2_G0_14_s0), .output_share1(d2_G0_14_s1));
  reg_module u_reg_G0_15_d2 (.clk(clk), .input_share0(d1_G0_15_s0), .input_share1(d1_G0_15_s1), .output_share0(d2_G0_15_s0), .output_share1(d2_G0_15_s1));
  reg_module u_reg_G0_16_d2 (.clk(clk), .input_share0(d1_G0_16_s0), .input_share1(d1_G0_16_s1), .output_share0(d2_G0_16_s0), .output_share1(d2_G0_16_s1));
  reg_module u_reg_G0_17_d2 (.clk(clk), .input_share0(d1_G0_17_s0), .input_share1(d1_G0_17_s1), .output_share0(d2_G0_17_s0), .output_share1(d2_G0_17_s1));
  reg_module u_reg_G0_18_d2 (.clk(clk), .input_share0(d1_G0_18_s0), .input_share1(d1_G0_18_s1), .output_share0(d2_G0_18_s0), .output_share1(d2_G0_18_s1));
  reg_module u_reg_G0_19_d2 (.clk(clk), .input_share0(d1_G0_19_s0), .input_share1(d1_G0_19_s1), .output_share0(d2_G0_19_s0), .output_share1(d2_G0_19_s1));
  reg_module u_reg_G0_2_d2 (.clk(clk), .input_share0(d1_G0_2_s0), .input_share1(d1_G0_2_s1), .output_share0(d2_G0_2_s0), .output_share1(d2_G0_2_s1));
  reg_module u_reg_G0_20_d2 (.clk(clk), .input_share0(d1_G0_20_s0), .input_share1(d1_G0_20_s1), .output_share0(d2_G0_20_s0), .output_share1(d2_G0_20_s1));
  reg_module u_reg_G0_21_d2 (.clk(clk), .input_share0(d1_G0_21_s0), .input_share1(d1_G0_21_s1), .output_share0(d2_G0_21_s0), .output_share1(d2_G0_21_s1));
  reg_module u_reg_G0_22_d2 (.clk(clk), .input_share0(d1_G0_22_s0), .input_share1(d1_G0_22_s1), .output_share0(d2_G0_22_s0), .output_share1(d2_G0_22_s1));
  reg_module u_reg_G0_23_d2 (.clk(clk), .input_share0(d1_G0_23_s0), .input_share1(d1_G0_23_s1), .output_share0(d2_G0_23_s0), .output_share1(d2_G0_23_s1));
  reg_module u_reg_G0_24_d2 (.clk(clk), .input_share0(d1_G0_24_s0), .input_share1(d1_G0_24_s1), .output_share0(d2_G0_24_s0), .output_share1(d2_G0_24_s1));
  reg_module u_reg_G0_25_d2 (.clk(clk), .input_share0(d1_G0_25_s0), .input_share1(d1_G0_25_s1), .output_share0(d2_G0_25_s0), .output_share1(d2_G0_25_s1));
  reg_module u_reg_G0_26_d2 (.clk(clk), .input_share0(d1_G0_26_s0), .input_share1(d1_G0_26_s1), .output_share0(d2_G0_26_s0), .output_share1(d2_G0_26_s1));
  reg_module u_reg_G0_27_d2 (.clk(clk), .input_share0(d1_G0_27_s0), .input_share1(d1_G0_27_s1), .output_share0(d2_G0_27_s0), .output_share1(d2_G0_27_s1));
  reg_module u_reg_G0_28_d2 (.clk(clk), .input_share0(d1_G0_28_s0), .input_share1(d1_G0_28_s1), .output_share0(d2_G0_28_s0), .output_share1(d2_G0_28_s1));
  reg_module u_reg_G0_29_d2 (.clk(clk), .input_share0(d1_G0_29_s0), .input_share1(d1_G0_29_s1), .output_share0(d2_G0_29_s0), .output_share1(d2_G0_29_s1));
  reg_module u_reg_G0_3_d2 (.clk(clk), .input_share0(d1_G0_3_s0), .input_share1(d1_G0_3_s1), .output_share0(d2_G0_3_s0), .output_share1(d2_G0_3_s1));
  reg_module u_reg_G0_30_d2 (.clk(clk), .input_share0(d1_G0_30_s0), .input_share1(d1_G0_30_s1), .output_share0(d2_G0_30_s0), .output_share1(d2_G0_30_s1));
  reg_module u_reg_G0_31_d2 (.clk(clk), .input_share0(d1_G0_31_s0), .input_share1(d1_G0_31_s1), .output_share0(d2_G0_31_s0), .output_share1(d2_G0_31_s1));
  reg_module u_reg_G0_4_d2 (.clk(clk), .input_share0(d1_G0_4_s0), .input_share1(d1_G0_4_s1), .output_share0(d2_G0_4_s0), .output_share1(d2_G0_4_s1));
  reg_module u_reg_G0_5_d2 (.clk(clk), .input_share0(d1_G0_5_s0), .input_share1(d1_G0_5_s1), .output_share0(d2_G0_5_s0), .output_share1(d2_G0_5_s1));
  reg_module u_reg_G0_6_d2 (.clk(clk), .input_share0(d1_G0_6_s0), .input_share1(d1_G0_6_s1), .output_share0(d2_G0_6_s0), .output_share1(d2_G0_6_s1));
  reg_module u_reg_G0_7_d2 (.clk(clk), .input_share0(d1_G0_7_s0), .input_share1(d1_G0_7_s1), .output_share0(d2_G0_7_s0), .output_share1(d2_G0_7_s1));
  reg_module u_reg_G0_8_d2 (.clk(clk), .input_share0(d1_G0_8_s0), .input_share1(d1_G0_8_s1), .output_share0(d2_G0_8_s0), .output_share1(d2_G0_8_s1));
  reg_module u_reg_G0_9_d2 (.clk(clk), .input_share0(d1_G0_9_s0), .input_share1(d1_G0_9_s1), .output_share0(d2_G0_9_s0), .output_share1(d2_G0_9_s1));
  reg_module u_reg_P0_10_d2 (.clk(clk), .input_share0(d1_P0_10_s0), .input_share1(d1_P0_10_s1), .output_share0(d2_P0_10_s0), .output_share1(d2_P0_10_s1));
  reg_module u_reg_P0_11_d2 (.clk(clk), .input_share0(d1_P0_11_s0), .input_share1(d1_P0_11_s1), .output_share0(d2_P0_11_s0), .output_share1(d2_P0_11_s1));
  reg_module u_reg_P0_12_d2 (.clk(clk), .input_share0(d1_P0_12_s0), .input_share1(d1_P0_12_s1), .output_share0(d2_P0_12_s0), .output_share1(d2_P0_12_s1));
  reg_module u_reg_P0_13_d2 (.clk(clk), .input_share0(d1_P0_13_s0), .input_share1(d1_P0_13_s1), .output_share0(d2_P0_13_s0), .output_share1(d2_P0_13_s1));
  reg_module u_reg_P0_14_d2 (.clk(clk), .input_share0(d1_P0_14_s0), .input_share1(d1_P0_14_s1), .output_share0(d2_P0_14_s0), .output_share1(d2_P0_14_s1));
  reg_module u_reg_P0_15_d2 (.clk(clk), .input_share0(d1_P0_15_s0), .input_share1(d1_P0_15_s1), .output_share0(d2_P0_15_s0), .output_share1(d2_P0_15_s1));
  reg_module u_reg_P0_16_d2 (.clk(clk), .input_share0(d1_P0_16_s0), .input_share1(d1_P0_16_s1), .output_share0(d2_P0_16_s0), .output_share1(d2_P0_16_s1));
  reg_module u_reg_P0_17_d2 (.clk(clk), .input_share0(d1_P0_17_s0), .input_share1(d1_P0_17_s1), .output_share0(d2_P0_17_s0), .output_share1(d2_P0_17_s1));
  reg_module u_reg_P0_18_d2 (.clk(clk), .input_share0(d1_P0_18_s0), .input_share1(d1_P0_18_s1), .output_share0(d2_P0_18_s0), .output_share1(d2_P0_18_s1));
  reg_module u_reg_P0_19_d2 (.clk(clk), .input_share0(d1_P0_19_s0), .input_share1(d1_P0_19_s1), .output_share0(d2_P0_19_s0), .output_share1(d2_P0_19_s1));
  reg_module u_reg_P0_2_d2 (.clk(clk), .input_share0(d1_P0_2_s0), .input_share1(d1_P0_2_s1), .output_share0(d2_P0_2_s0), .output_share1(d2_P0_2_s1));
  reg_module u_reg_P0_20_d2 (.clk(clk), .input_share0(d1_P0_20_s0), .input_share1(d1_P0_20_s1), .output_share0(d2_P0_20_s0), .output_share1(d2_P0_20_s1));
  reg_module u_reg_P0_21_d2 (.clk(clk), .input_share0(d1_P0_21_s0), .input_share1(d1_P0_21_s1), .output_share0(d2_P0_21_s0), .output_share1(d2_P0_21_s1));
  reg_module u_reg_P0_22_d2 (.clk(clk), .input_share0(d1_P0_22_s0), .input_share1(d1_P0_22_s1), .output_share0(d2_P0_22_s0), .output_share1(d2_P0_22_s1));
  reg_module u_reg_P0_23_d2 (.clk(clk), .input_share0(d1_P0_23_s0), .input_share1(d1_P0_23_s1), .output_share0(d2_P0_23_s0), .output_share1(d2_P0_23_s1));
  reg_module u_reg_P0_24_d2 (.clk(clk), .input_share0(d1_P0_24_s0), .input_share1(d1_P0_24_s1), .output_share0(d2_P0_24_s0), .output_share1(d2_P0_24_s1));
  reg_module u_reg_P0_25_d2 (.clk(clk), .input_share0(d1_P0_25_s0), .input_share1(d1_P0_25_s1), .output_share0(d2_P0_25_s0), .output_share1(d2_P0_25_s1));
  reg_module u_reg_P0_26_d2 (.clk(clk), .input_share0(d1_P0_26_s0), .input_share1(d1_P0_26_s1), .output_share0(d2_P0_26_s0), .output_share1(d2_P0_26_s1));
  reg_module u_reg_P0_27_d2 (.clk(clk), .input_share0(d1_P0_27_s0), .input_share1(d1_P0_27_s1), .output_share0(d2_P0_27_s0), .output_share1(d2_P0_27_s1));
  reg_module u_reg_P0_28_d2 (.clk(clk), .input_share0(d1_P0_28_s0), .input_share1(d1_P0_28_s1), .output_share0(d2_P0_28_s0), .output_share1(d2_P0_28_s1));
  reg_module u_reg_P0_29_d2 (.clk(clk), .input_share0(d1_P0_29_s0), .input_share1(d1_P0_29_s1), .output_share0(d2_P0_29_s0), .output_share1(d2_P0_29_s1));
  reg_module u_reg_P0_3_d2 (.clk(clk), .input_share0(d1_P0_3_s0), .input_share1(d1_P0_3_s1), .output_share0(d2_P0_3_s0), .output_share1(d2_P0_3_s1));
  reg_module u_reg_P0_30_d2 (.clk(clk), .input_share0(d1_P0_30_s0), .input_share1(d1_P0_30_s1), .output_share0(d2_P0_30_s0), .output_share1(d2_P0_30_s1));
  reg_module u_reg_P0_31_d2 (.clk(clk), .input_share0(d1_P0_31_s0), .input_share1(d1_P0_31_s1), .output_share0(d2_P0_31_s0), .output_share1(d2_P0_31_s1));
  reg_module u_reg_P0_4_d2 (.clk(clk), .input_share0(d1_P0_4_s0), .input_share1(d1_P0_4_s1), .output_share0(d2_P0_4_s0), .output_share1(d2_P0_4_s1));
  reg_module u_reg_P0_5_d2 (.clk(clk), .input_share0(d1_P0_5_s0), .input_share1(d1_P0_5_s1), .output_share0(d2_P0_5_s0), .output_share1(d2_P0_5_s1));
  reg_module u_reg_P0_6_d2 (.clk(clk), .input_share0(d1_P0_6_s0), .input_share1(d1_P0_6_s1), .output_share0(d2_P0_6_s0), .output_share1(d2_P0_6_s1));
  reg_module u_reg_P0_7_d2 (.clk(clk), .input_share0(d1_P0_7_s0), .input_share1(d1_P0_7_s1), .output_share0(d2_P0_7_s0), .output_share1(d2_P0_7_s1));
  reg_module u_reg_P0_8_d2 (.clk(clk), .input_share0(d1_P0_8_s0), .input_share1(d1_P0_8_s1), .output_share0(d2_P0_8_s0), .output_share1(d2_P0_8_s1));
  reg_module u_reg_P0_9_d2 (.clk(clk), .input_share0(d1_P0_9_s0), .input_share1(d1_P0_9_s1), .output_share0(d2_P0_9_s0), .output_share1(d2_P0_9_s1));
  reg_module u_reg_P1_11_d2 (.clk(clk), .input_share0(d1_P1_11_s0), .input_share1(d1_P1_11_s1), .output_share0(d2_P1_11_s0), .output_share1(d2_P1_11_s1));
  reg_module u_reg_P1_13_d2 (.clk(clk), .input_share0(d1_P1_13_s0), .input_share1(d1_P1_13_s1), .output_share0(d2_P1_13_s0), .output_share1(d2_P1_13_s1));
  reg_module u_reg_P1_15_d2 (.clk(clk), .input_share0(d1_P1_15_s0), .input_share1(d1_P1_15_s1), .output_share0(d2_P1_15_s0), .output_share1(d2_P1_15_s1));
  reg_module u_reg_P1_17_d2 (.clk(clk), .input_share0(d1_P1_17_s0), .input_share1(d1_P1_17_s1), .output_share0(d2_P1_17_s0), .output_share1(d2_P1_17_s1));
  reg_module u_reg_P1_19_d2 (.clk(clk), .input_share0(d1_P1_19_s0), .input_share1(d1_P1_19_s1), .output_share0(d2_P1_19_s0), .output_share1(d2_P1_19_s1));
  reg_module u_reg_P1_21_d2 (.clk(clk), .input_share0(d1_P1_21_s0), .input_share1(d1_P1_21_s1), .output_share0(d2_P1_21_s0), .output_share1(d2_P1_21_s1));
  reg_module u_reg_P1_23_d2 (.clk(clk), .input_share0(d1_P1_23_s0), .input_share1(d1_P1_23_s1), .output_share0(d2_P1_23_s0), .output_share1(d2_P1_23_s1));
  reg_module u_reg_P1_25_d2 (.clk(clk), .input_share0(d1_P1_25_s0), .input_share1(d1_P1_25_s1), .output_share0(d2_P1_25_s0), .output_share1(d2_P1_25_s1));
  reg_module u_reg_P1_27_d2 (.clk(clk), .input_share0(d1_P1_27_s0), .input_share1(d1_P1_27_s1), .output_share0(d2_P1_27_s0), .output_share1(d2_P1_27_s1));
  reg_module u_reg_P1_29_d2 (.clk(clk), .input_share0(d1_P1_29_s0), .input_share1(d1_P1_29_s1), .output_share0(d2_P1_29_s0), .output_share1(d2_P1_29_s1));
  reg_module u_reg_P1_3_d2 (.clk(clk), .input_share0(d1_P1_3_s0), .input_share1(d1_P1_3_s1), .output_share0(d2_P1_3_s0), .output_share1(d2_P1_3_s1));
  reg_module u_reg_P1_31_d2 (.clk(clk), .input_share0(d1_P1_31_s0), .input_share1(d1_P1_31_s1), .output_share0(d2_P1_31_s0), .output_share1(d2_P1_31_s1));
  reg_module u_reg_P1_5_d2 (.clk(clk), .input_share0(d1_P1_5_s0), .input_share1(d1_P1_5_s1), .output_share0(d2_P1_5_s0), .output_share1(d2_P1_5_s1));
  reg_module u_reg_P1_7_d2 (.clk(clk), .input_share0(d1_P1_7_s0), .input_share1(d1_P1_7_s1), .output_share0(d2_P1_7_s0), .output_share1(d2_P1_7_s1));
  reg_module u_reg_P1_9_d2 (.clk(clk), .input_share0(d1_P1_9_s0), .input_share1(d1_P1_9_s1), .output_share0(d2_P1_9_s0), .output_share1(d2_P1_9_s1));
  xor_module u_xor_G1_1_d2 (.x_share0(d2_t0_s0), .x_share1(d2_t0_s1), .y_share0(d2_G0_1_s0), .y_share1(d2_G0_1_s1), .z_share0(d2_G1_1_s0), .z_share1(d2_G1_1_s1));
  xor_module u_xor_G1_11_d2 (.x_share0(d2_t5_s0), .x_share1(d2_t5_s1), .y_share0(d2_G0_11_s0), .y_share1(d2_G0_11_s1), .z_share0(d2_G1_11_s0), .z_share1(d2_G1_11_s1));
  xor_module u_xor_G1_13_d2 (.x_share0(d2_t6_s0), .x_share1(d2_t6_s1), .y_share0(d2_G0_13_s0), .y_share1(d2_G0_13_s1), .z_share0(d2_G1_13_s0), .z_share1(d2_G1_13_s1));
  xor_module u_xor_G1_15_d2 (.x_share0(d2_t7_s0), .x_share1(d2_t7_s1), .y_share0(d2_G0_15_s0), .y_share1(d2_G0_15_s1), .z_share0(d2_G1_15_s0), .z_share1(d2_G1_15_s1));
  xor_module u_xor_G1_17_d2 (.x_share0(d2_t8_s0), .x_share1(d2_t8_s1), .y_share0(d2_G0_17_s0), .y_share1(d2_G0_17_s1), .z_share0(d2_G1_17_s0), .z_share1(d2_G1_17_s1));
  xor_module u_xor_G1_19_d2 (.x_share0(d2_t9_s0), .x_share1(d2_t9_s1), .y_share0(d2_G0_19_s0), .y_share1(d2_G0_19_s1), .z_share0(d2_G1_19_s0), .z_share1(d2_G1_19_s1));
  xor_module u_xor_G1_21_d2 (.x_share0(d2_t10_s0), .x_share1(d2_t10_s1), .y_share0(d2_G0_21_s0), .y_share1(d2_G0_21_s1), .z_share0(d2_G1_21_s0), .z_share1(d2_G1_21_s1));
  xor_module u_xor_G1_23_d2 (.x_share0(d2_t11_s0), .x_share1(d2_t11_s1), .y_share0(d2_G0_23_s0), .y_share1(d2_G0_23_s1), .z_share0(d2_G1_23_s0), .z_share1(d2_G1_23_s1));
  xor_module u_xor_G1_25_d2 (.x_share0(d2_t12_s0), .x_share1(d2_t12_s1), .y_share0(d2_G0_25_s0), .y_share1(d2_G0_25_s1), .z_share0(d2_G1_25_s0), .z_share1(d2_G1_25_s1));
  xor_module u_xor_G1_27_d2 (.x_share0(d2_t13_s0), .x_share1(d2_t13_s1), .y_share0(d2_G0_27_s0), .y_share1(d2_G0_27_s1), .z_share0(d2_G1_27_s0), .z_share1(d2_G1_27_s1));
  xor_module u_xor_G1_29_d2 (.x_share0(d2_t14_s0), .x_share1(d2_t14_s1), .y_share0(d2_G0_29_s0), .y_share1(d2_G0_29_s1), .z_share0(d2_G1_29_s0), .z_share1(d2_G1_29_s1));
  xor_module u_xor_G1_3_d2 (.x_share0(d2_t1_s0), .x_share1(d2_t1_s1), .y_share0(d2_G0_3_s0), .y_share1(d2_G0_3_s1), .z_share0(d2_G1_3_s0), .z_share1(d2_G1_3_s1));
  xor_module u_xor_G1_31_d2 (.x_share0(d2_t15_s0), .x_share1(d2_t15_s1), .y_share0(d2_G0_31_s0), .y_share1(d2_G0_31_s1), .z_share0(d2_G1_31_s0), .z_share1(d2_G1_31_s1));
  xor_module u_xor_G1_5_d2 (.x_share0(d2_t2_s0), .x_share1(d2_t2_s1), .y_share0(d2_G0_5_s0), .y_share1(d2_G0_5_s1), .z_share0(d2_G1_5_s0), .z_share1(d2_G1_5_s1));
  xor_module u_xor_G1_7_d2 (.x_share0(d2_t3_s0), .x_share1(d2_t3_s1), .y_share0(d2_G0_7_s0), .y_share1(d2_G0_7_s1), .z_share0(d2_G1_7_s0), .z_share1(d2_G1_7_s1));
  xor_module u_xor_G1_9_d2 (.x_share0(d2_t4_s0), .x_share1(d2_t4_s1), .y_share0(d2_G0_9_s0), .y_share1(d2_G0_9_s1), .z_share0(d2_G1_9_s0), .z_share1(d2_G1_9_s1));
  and_module u_and_P2_10_d2 (.clk(clk), .x_share0(d1_P0_10_s0), .x_share1(d1_P0_10_s1), .y_share0(d1_P1_9_s0), .y_share1(d1_P1_9_s1), .rand(r_P2_10), .z_share0(d2_P2_10_s0), .z_share1(d2_P2_10_s1));
  assign r_P2_10 = stage2_share0[0];
  and_module u_and_P2_11_d2 (.clk(clk), .x_share0(d1_P1_11_s0), .x_share1(d1_P1_11_s1), .y_share0(d1_P1_9_s0), .y_share1(d1_P1_9_s1), .rand(r_P2_11), .z_share0(d2_P2_11_s0), .z_share1(d2_P2_11_s1));
  assign r_P2_11 = stage2_share0[4];
  and_module u_and_P2_14_d2 (.clk(clk), .x_share0(d1_P0_14_s0), .x_share1(d1_P0_14_s1), .y_share0(d1_P1_13_s0), .y_share1(d1_P1_13_s1), .rand(r_P2_14), .z_share0(d2_P2_14_s0), .z_share1(d2_P2_14_s1));
  assign r_P2_14 = stage2_share0[1];
  and_module u_and_P2_15_d2 (.clk(clk), .x_share0(d1_P1_15_s0), .x_share1(d1_P1_15_s1), .y_share0(d1_P1_13_s0), .y_share1(d1_P1_13_s1), .rand(r_P2_15), .z_share0(d2_P2_15_s0), .z_share1(d2_P2_15_s1));
  assign r_P2_15 = stage2_share0[1];
  and_module u_and_P2_18_d2 (.clk(clk), .x_share0(d1_P0_18_s0), .x_share1(d1_P0_18_s1), .y_share0(d1_P1_17_s0), .y_share1(d1_P1_17_s1), .rand(r_P2_18), .z_share0(d2_P2_18_s0), .z_share1(d2_P2_18_s1));
  assign r_P2_18 = stage2_share0[14];
  and_module u_and_P2_19_d2 (.clk(clk), .x_share0(d1_P1_19_s0), .x_share1(d1_P1_19_s1), .y_share0(d1_P1_17_s0), .y_share1(d1_P1_17_s1), .rand(r_P2_19), .z_share0(d2_P2_19_s0), .z_share1(d2_P2_19_s1));
  assign r_P2_19 = stage2_share0[18];
  and_module u_and_P2_22_d2 (.clk(clk), .x_share0(d1_P0_22_s0), .x_share1(d1_P0_22_s1), .y_share0(d1_P1_21_s0), .y_share1(d1_P1_21_s1), .rand(r_P2_22), .z_share0(d2_P2_22_s0), .z_share1(d2_P2_22_s1));
  assign r_P2_22 = stage2_share0[14];
  and_module u_and_P2_23_d2 (.clk(clk), .x_share0(d1_P1_23_s0), .x_share1(d1_P1_23_s1), .y_share0(d1_P1_21_s0), .y_share1(d1_P1_21_s1), .rand(r_P2_23), .z_share0(d2_P2_23_s0), .z_share1(d2_P2_23_s1));
  assign r_P2_23 = stage2_share0[15];
  and_module u_and_P2_26_d2 (.clk(clk), .x_share0(d1_P0_26_s0), .x_share1(d1_P0_26_s1), .y_share0(d1_P1_25_s0), .y_share1(d1_P1_25_s1), .rand(r_P2_26), .z_share0(d2_P2_26_s0), .z_share1(d2_P2_26_s1));
  assign r_P2_26 = stage2_share0[17];
  and_module u_and_P2_27_d2 (.clk(clk), .x_share0(d1_P1_27_s0), .x_share1(d1_P1_27_s1), .y_share0(d1_P1_25_s0), .y_share1(d1_P1_25_s1), .rand(r_P2_27), .z_share0(d2_P2_27_s0), .z_share1(d2_P2_27_s1));
  assign r_P2_27 = stage2_share0[21];
  and_module u_and_P2_30_d2 (.clk(clk), .x_share0(d1_P0_30_s0), .x_share1(d1_P0_30_s1), .y_share0(d1_P1_29_s0), .y_share1(d1_P1_29_s1), .rand(r_P2_30), .z_share0(d2_P2_30_s0), .z_share1(d2_P2_30_s1));
  assign r_P2_30 = stage2_share0[19];
  and_module u_and_P2_31_d2 (.clk(clk), .x_share0(d1_P1_31_s0), .x_share1(d1_P1_31_s1), .y_share0(d1_P1_29_s0), .y_share1(d1_P1_29_s1), .rand(r_P2_31), .z_share0(d2_P2_31_s0), .z_share1(d2_P2_31_s1));
  assign r_P2_31 = stage2_share0[23];
  and_module u_and_P2_6_d2 (.clk(clk), .x_share0(d1_P0_6_s0), .x_share1(d1_P0_6_s1), .y_share0(d1_P1_5_s0), .y_share1(d1_P1_5_s1), .rand(r_P2_6), .z_share0(d2_P2_6_s0), .z_share1(d2_P2_6_s1));
  assign r_P2_6 = stage2_share0[3];
  and_module u_and_P2_7_d2 (.clk(clk), .x_share0(d1_P1_7_s0), .x_share1(d1_P1_7_s1), .y_share0(d1_P1_5_s0), .y_share1(d1_P1_5_s1), .rand(r_P2_7), .z_share0(d2_P2_7_s0), .z_share1(d2_P2_7_s1));
  assign r_P2_7 = stage2_share0[10];
  xor_module u_xor_o2_d2 (.x_share0(d2_P0_2_s0), .x_share1(d2_P0_2_s1), .y_share0(d2_G1_1_s0), .y_share1(d2_G1_1_s1), .z_share0(d2_o2_s0), .z_share1(d2_o2_s1));
  and_module u_and_t0_d2 (.clk(clk), .x_share0(d1_P0_1_s0), .x_share1(d1_P0_1_s1), .y_share0(d1_G0_0_s0), .y_share1(d1_G0_0_s1), .rand(r_t0), .z_share0(d2_t0_s0), .z_share1(d2_t0_s1));
  assign r_t0 = stage2_share0[1];
  and_module u_and_t1_d2 (.clk(clk), .x_share0(d1_P0_3_s0), .x_share1(d1_P0_3_s1), .y_share0(d1_G0_2_s0), .y_share1(d1_G0_2_s1), .rand(r_t1), .z_share0(d2_t1_s0), .z_share1(d2_t1_s1));
  assign r_t1 = stage2_share0[15];
  and_module u_and_t10_d2 (.clk(clk), .x_share0(d1_P0_21_s0), .x_share1(d1_P0_21_s1), .y_share0(d1_G0_20_s0), .y_share1(d1_G0_20_s1), .rand(r_t10), .z_share0(d2_t10_s0), .z_share1(d2_t10_s1));
  assign r_t10 = stage2_share0[15];
  and_module u_and_t11_d2 (.clk(clk), .x_share0(d1_P0_23_s0), .x_share1(d1_P0_23_s1), .y_share0(d1_G0_22_s0), .y_share1(d1_G0_22_s1), .rand(r_t11), .z_share0(d2_t11_s0), .z_share1(d2_t11_s1));
  assign r_t11 = stage2_share0[9];
  and_module u_and_t12_d2 (.clk(clk), .x_share0(d1_P0_25_s0), .x_share1(d1_P0_25_s1), .y_share0(d1_G0_24_s0), .y_share1(d1_G0_24_s1), .rand(r_t12), .z_share0(d2_t12_s0), .z_share1(d2_t12_s1));
  assign r_t12 = stage2_share0[21];
  and_module u_and_t13_d2 (.clk(clk), .x_share0(d1_P0_27_s0), .x_share1(d1_P0_27_s1), .y_share0(d1_G0_26_s0), .y_share1(d1_G0_26_s1), .rand(r_t13), .z_share0(d2_t13_s0), .z_share1(d2_t13_s1));
  assign r_t13 = stage2_share0[13];
  and_module u_and_t14_d2 (.clk(clk), .x_share0(d1_P0_29_s0), .x_share1(d1_P0_29_s1), .y_share0(d1_G0_28_s0), .y_share1(d1_G0_28_s1), .rand(r_t14), .z_share0(d2_t14_s0), .z_share1(d2_t14_s1));
  assign r_t14 = stage2_share0[25];
  and_module u_and_t15_d2 (.clk(clk), .x_share0(d1_P0_31_s0), .x_share1(d1_P0_31_s1), .y_share0(d1_G0_30_s0), .y_share1(d1_G0_30_s1), .rand(r_t15), .z_share0(d2_t15_s0), .z_share1(d2_t15_s1));
  assign r_t15 = stage2_share0[21];
  and_module u_and_t2_d2 (.clk(clk), .x_share0(d1_P0_5_s0), .x_share1(d1_P0_5_s1), .y_share0(d1_G0_4_s0), .y_share1(d1_G0_4_s1), .rand(r_t2), .z_share0(d2_t2_s0), .z_share1(d2_t2_s1));
  assign r_t2 = stage2_share0[1];
  and_module u_and_t3_d2 (.clk(clk), .x_share0(d1_P0_7_s0), .x_share1(d1_P0_7_s1), .y_share0(d1_G0_6_s0), .y_share1(d1_G0_6_s1), .rand(r_t3), .z_share0(d2_t3_s0), .z_share1(d2_t3_s1));
  assign r_t3 = stage2_share0[11];
  and_module u_and_t4_d2 (.clk(clk), .x_share0(d1_P0_9_s0), .x_share1(d1_P0_9_s1), .y_share0(d1_G0_8_s0), .y_share1(d1_G0_8_s1), .rand(r_t4), .z_share0(d2_t4_s0), .z_share1(d2_t4_s1));
  assign r_t4 = stage2_share0[5];
  and_module u_and_t5_d2 (.clk(clk), .x_share0(d1_P0_11_s0), .x_share1(d1_P0_11_s1), .y_share0(d1_G0_10_s0), .y_share1(d1_G0_10_s1), .rand(r_t5), .z_share0(d2_t5_s0), .z_share1(d2_t5_s1));
  assign r_t5 = stage2_share0[14];
  and_module u_and_t6_d2 (.clk(clk), .x_share0(d1_P0_13_s0), .x_share1(d1_P0_13_s1), .y_share0(d1_G0_12_s0), .y_share1(d1_G0_12_s1), .rand(r_t6), .z_share0(d2_t6_s0), .z_share1(d2_t6_s1));
  assign r_t6 = stage2_share0[6];
  and_module u_and_t7_d2 (.clk(clk), .x_share0(d1_P0_15_s0), .x_share1(d1_P0_15_s1), .y_share0(d1_G0_14_s0), .y_share1(d1_G0_14_s1), .rand(r_t7), .z_share0(d2_t7_s0), .z_share1(d2_t7_s1));
  assign r_t7 = stage2_share0[4];
  and_module u_and_t8_d2 (.clk(clk), .x_share0(d1_P0_17_s0), .x_share1(d1_P0_17_s1), .y_share0(d1_G0_16_s0), .y_share1(d1_G0_16_s1), .rand(r_t8), .z_share0(d2_t8_s0), .z_share1(d2_t8_s1));
  assign r_t8 = stage2_share0[9];
  and_module u_and_t9_d2 (.clk(clk), .x_share0(d1_P0_19_s0), .x_share1(d1_P0_19_s1), .y_share0(d1_G0_18_s0), .y_share1(d1_G0_18_s1), .rand(r_t9), .z_share0(d2_t9_s0), .z_share1(d2_t9_s1));
  assign r_t9 = stage2_share0[13];
  reg_module u_reg_G0_10_d3 (.clk(clk), .input_share0(d2_G0_10_s0), .input_share1(d2_G0_10_s1), .output_share0(d3_G0_10_s0), .output_share1(d3_G0_10_s1));
  reg_module u_reg_G0_12_d3 (.clk(clk), .input_share0(d2_G0_12_s0), .input_share1(d2_G0_12_s1), .output_share0(d3_G0_12_s0), .output_share1(d3_G0_12_s1));
  reg_module u_reg_G0_14_d3 (.clk(clk), .input_share0(d2_G0_14_s0), .input_share1(d2_G0_14_s1), .output_share0(d3_G0_14_s0), .output_share1(d3_G0_14_s1));
  reg_module u_reg_G0_16_d3 (.clk(clk), .input_share0(d2_G0_16_s0), .input_share1(d2_G0_16_s1), .output_share0(d3_G0_16_s0), .output_share1(d3_G0_16_s1));
  reg_module u_reg_G0_18_d3 (.clk(clk), .input_share0(d2_G0_18_s0), .input_share1(d2_G0_18_s1), .output_share0(d3_G0_18_s0), .output_share1(d3_G0_18_s1));
  reg_module u_reg_G0_2_d3 (.clk(clk), .input_share0(d2_G0_2_s0), .input_share1(d2_G0_2_s1), .output_share0(d3_G0_2_s0), .output_share1(d3_G0_2_s1));
  reg_module u_reg_G0_20_d3 (.clk(clk), .input_share0(d2_G0_20_s0), .input_share1(d2_G0_20_s1), .output_share0(d3_G0_20_s0), .output_share1(d3_G0_20_s1));
  reg_module u_reg_G0_22_d3 (.clk(clk), .input_share0(d2_G0_22_s0), .input_share1(d2_G0_22_s1), .output_share0(d3_G0_22_s0), .output_share1(d3_G0_22_s1));
  reg_module u_reg_G0_24_d3 (.clk(clk), .input_share0(d2_G0_24_s0), .input_share1(d2_G0_24_s1), .output_share0(d3_G0_24_s0), .output_share1(d3_G0_24_s1));
  reg_module u_reg_G0_26_d3 (.clk(clk), .input_share0(d2_G0_26_s0), .input_share1(d2_G0_26_s1), .output_share0(d3_G0_26_s0), .output_share1(d3_G0_26_s1));
  reg_module u_reg_G0_28_d3 (.clk(clk), .input_share0(d2_G0_28_s0), .input_share1(d2_G0_28_s1), .output_share0(d3_G0_28_s0), .output_share1(d3_G0_28_s1));
  reg_module u_reg_G0_30_d3 (.clk(clk), .input_share0(d2_G0_30_s0), .input_share1(d2_G0_30_s1), .output_share0(d3_G0_30_s0), .output_share1(d3_G0_30_s1));
  reg_module u_reg_G0_4_d3 (.clk(clk), .input_share0(d2_G0_4_s0), .input_share1(d2_G0_4_s1), .output_share0(d3_G0_4_s0), .output_share1(d3_G0_4_s1));
  reg_module u_reg_G0_6_d3 (.clk(clk), .input_share0(d2_G0_6_s0), .input_share1(d2_G0_6_s1), .output_share0(d3_G0_6_s0), .output_share1(d3_G0_6_s1));
  reg_module u_reg_G0_8_d3 (.clk(clk), .input_share0(d2_G0_8_s0), .input_share1(d2_G0_8_s1), .output_share0(d3_G0_8_s0), .output_share1(d3_G0_8_s1));
  reg_module u_reg_G1_11_d3 (.clk(clk), .input_share0(d2_G1_11_s0), .input_share1(d2_G1_11_s1), .output_share0(d3_G1_11_s0), .output_share1(d3_G1_11_s1));
  reg_module u_reg_G1_13_d3 (.clk(clk), .input_share0(d2_G1_13_s0), .input_share1(d2_G1_13_s1), .output_share0(d3_G1_13_s0), .output_share1(d3_G1_13_s1));
  reg_module u_reg_G1_15_d3 (.clk(clk), .input_share0(d2_G1_15_s0), .input_share1(d2_G1_15_s1), .output_share0(d3_G1_15_s0), .output_share1(d3_G1_15_s1));
  reg_module u_reg_G1_17_d3 (.clk(clk), .input_share0(d2_G1_17_s0), .input_share1(d2_G1_17_s1), .output_share0(d3_G1_17_s0), .output_share1(d3_G1_17_s1));
  reg_module u_reg_G1_19_d3 (.clk(clk), .input_share0(d2_G1_19_s0), .input_share1(d2_G1_19_s1), .output_share0(d3_G1_19_s0), .output_share1(d3_G1_19_s1));
  reg_module u_reg_G1_21_d3 (.clk(clk), .input_share0(d2_G1_21_s0), .input_share1(d2_G1_21_s1), .output_share0(d3_G1_21_s0), .output_share1(d3_G1_21_s1));
  reg_module u_reg_G1_23_d3 (.clk(clk), .input_share0(d2_G1_23_s0), .input_share1(d2_G1_23_s1), .output_share0(d3_G1_23_s0), .output_share1(d3_G1_23_s1));
  reg_module u_reg_G1_25_d3 (.clk(clk), .input_share0(d2_G1_25_s0), .input_share1(d2_G1_25_s1), .output_share0(d3_G1_25_s0), .output_share1(d3_G1_25_s1));
  reg_module u_reg_G1_27_d3 (.clk(clk), .input_share0(d2_G1_27_s0), .input_share1(d2_G1_27_s1), .output_share0(d3_G1_27_s0), .output_share1(d3_G1_27_s1));
  reg_module u_reg_G1_29_d3 (.clk(clk), .input_share0(d2_G1_29_s0), .input_share1(d2_G1_29_s1), .output_share0(d3_G1_29_s0), .output_share1(d3_G1_29_s1));
  reg_module u_reg_G1_3_d3 (.clk(clk), .input_share0(d2_G1_3_s0), .input_share1(d2_G1_3_s1), .output_share0(d3_G1_3_s0), .output_share1(d3_G1_3_s1));
  reg_module u_reg_G1_31_d3 (.clk(clk), .input_share0(d2_G1_31_s0), .input_share1(d2_G1_31_s1), .output_share0(d3_G1_31_s0), .output_share1(d3_G1_31_s1));
  reg_module u_reg_G1_5_d3 (.clk(clk), .input_share0(d2_G1_5_s0), .input_share1(d2_G1_5_s1), .output_share0(d3_G1_5_s0), .output_share1(d3_G1_5_s1));
  reg_module u_reg_G1_7_d3 (.clk(clk), .input_share0(d2_G1_7_s0), .input_share1(d2_G1_7_s1), .output_share0(d3_G1_7_s0), .output_share1(d3_G1_7_s1));
  reg_module u_reg_G1_9_d3 (.clk(clk), .input_share0(d2_G1_9_s0), .input_share1(d2_G1_9_s1), .output_share0(d3_G1_9_s0), .output_share1(d3_G1_9_s1));
  reg_module u_reg_P0_10_d3 (.clk(clk), .input_share0(d2_P0_10_s0), .input_share1(d2_P0_10_s1), .output_share0(d3_P0_10_s0), .output_share1(d3_P0_10_s1));
  reg_module u_reg_P0_11_d3 (.clk(clk), .input_share0(d2_P0_11_s0), .input_share1(d2_P0_11_s1), .output_share0(d3_P0_11_s0), .output_share1(d3_P0_11_s1));
  reg_module u_reg_P0_12_d3 (.clk(clk), .input_share0(d2_P0_12_s0), .input_share1(d2_P0_12_s1), .output_share0(d3_P0_12_s0), .output_share1(d3_P0_12_s1));
  reg_module u_reg_P0_13_d3 (.clk(clk), .input_share0(d2_P0_13_s0), .input_share1(d2_P0_13_s1), .output_share0(d3_P0_13_s0), .output_share1(d3_P0_13_s1));
  reg_module u_reg_P0_14_d3 (.clk(clk), .input_share0(d2_P0_14_s0), .input_share1(d2_P0_14_s1), .output_share0(d3_P0_14_s0), .output_share1(d3_P0_14_s1));
  reg_module u_reg_P0_15_d3 (.clk(clk), .input_share0(d2_P0_15_s0), .input_share1(d2_P0_15_s1), .output_share0(d3_P0_15_s0), .output_share1(d3_P0_15_s1));
  reg_module u_reg_P0_16_d3 (.clk(clk), .input_share0(d2_P0_16_s0), .input_share1(d2_P0_16_s1), .output_share0(d3_P0_16_s0), .output_share1(d3_P0_16_s1));
  reg_module u_reg_P0_17_d3 (.clk(clk), .input_share0(d2_P0_17_s0), .input_share1(d2_P0_17_s1), .output_share0(d3_P0_17_s0), .output_share1(d3_P0_17_s1));
  reg_module u_reg_P0_18_d3 (.clk(clk), .input_share0(d2_P0_18_s0), .input_share1(d2_P0_18_s1), .output_share0(d3_P0_18_s0), .output_share1(d3_P0_18_s1));
  reg_module u_reg_P0_19_d3 (.clk(clk), .input_share0(d2_P0_19_s0), .input_share1(d2_P0_19_s1), .output_share0(d3_P0_19_s0), .output_share1(d3_P0_19_s1));
  reg_module u_reg_P0_20_d3 (.clk(clk), .input_share0(d2_P0_20_s0), .input_share1(d2_P0_20_s1), .output_share0(d3_P0_20_s0), .output_share1(d3_P0_20_s1));
  reg_module u_reg_P0_21_d3 (.clk(clk), .input_share0(d2_P0_21_s0), .input_share1(d2_P0_21_s1), .output_share0(d3_P0_21_s0), .output_share1(d3_P0_21_s1));
  reg_module u_reg_P0_22_d3 (.clk(clk), .input_share0(d2_P0_22_s0), .input_share1(d2_P0_22_s1), .output_share0(d3_P0_22_s0), .output_share1(d3_P0_22_s1));
  reg_module u_reg_P0_23_d3 (.clk(clk), .input_share0(d2_P0_23_s0), .input_share1(d2_P0_23_s1), .output_share0(d3_P0_23_s0), .output_share1(d3_P0_23_s1));
  reg_module u_reg_P0_24_d3 (.clk(clk), .input_share0(d2_P0_24_s0), .input_share1(d2_P0_24_s1), .output_share0(d3_P0_24_s0), .output_share1(d3_P0_24_s1));
  reg_module u_reg_P0_25_d3 (.clk(clk), .input_share0(d2_P0_25_s0), .input_share1(d2_P0_25_s1), .output_share0(d3_P0_25_s0), .output_share1(d3_P0_25_s1));
  reg_module u_reg_P0_26_d3 (.clk(clk), .input_share0(d2_P0_26_s0), .input_share1(d2_P0_26_s1), .output_share0(d3_P0_26_s0), .output_share1(d3_P0_26_s1));
  reg_module u_reg_P0_27_d3 (.clk(clk), .input_share0(d2_P0_27_s0), .input_share1(d2_P0_27_s1), .output_share0(d3_P0_27_s0), .output_share1(d3_P0_27_s1));
  reg_module u_reg_P0_28_d3 (.clk(clk), .input_share0(d2_P0_28_s0), .input_share1(d2_P0_28_s1), .output_share0(d3_P0_28_s0), .output_share1(d3_P0_28_s1));
  reg_module u_reg_P0_29_d3 (.clk(clk), .input_share0(d2_P0_29_s0), .input_share1(d2_P0_29_s1), .output_share0(d3_P0_29_s0), .output_share1(d3_P0_29_s1));
  reg_module u_reg_P0_3_d3 (.clk(clk), .input_share0(d2_P0_3_s0), .input_share1(d2_P0_3_s1), .output_share0(d3_P0_3_s0), .output_share1(d3_P0_3_s1));
  reg_module u_reg_P0_30_d3 (.clk(clk), .input_share0(d2_P0_30_s0), .input_share1(d2_P0_30_s1), .output_share0(d3_P0_30_s0), .output_share1(d3_P0_30_s1));
  reg_module u_reg_P0_31_d3 (.clk(clk), .input_share0(d2_P0_31_s0), .input_share1(d2_P0_31_s1), .output_share0(d3_P0_31_s0), .output_share1(d3_P0_31_s1));
  reg_module u_reg_P0_4_d3 (.clk(clk), .input_share0(d2_P0_4_s0), .input_share1(d2_P0_4_s1), .output_share0(d3_P0_4_s0), .output_share1(d3_P0_4_s1));
  reg_module u_reg_P0_5_d3 (.clk(clk), .input_share0(d2_P0_5_s0), .input_share1(d2_P0_5_s1), .output_share0(d3_P0_5_s0), .output_share1(d3_P0_5_s1));
  reg_module u_reg_P0_6_d3 (.clk(clk), .input_share0(d2_P0_6_s0), .input_share1(d2_P0_6_s1), .output_share0(d3_P0_6_s0), .output_share1(d3_P0_6_s1));
  reg_module u_reg_P0_7_d3 (.clk(clk), .input_share0(d2_P0_7_s0), .input_share1(d2_P0_7_s1), .output_share0(d3_P0_7_s0), .output_share1(d3_P0_7_s1));
  reg_module u_reg_P0_8_d3 (.clk(clk), .input_share0(d2_P0_8_s0), .input_share1(d2_P0_8_s1), .output_share0(d3_P0_8_s0), .output_share1(d3_P0_8_s1));
  reg_module u_reg_P0_9_d3 (.clk(clk), .input_share0(d2_P0_9_s0), .input_share1(d2_P0_9_s1), .output_share0(d3_P0_9_s0), .output_share1(d3_P0_9_s1));
  reg_module u_reg_P1_13_d3 (.clk(clk), .input_share0(d2_P1_13_s0), .input_share1(d2_P1_13_s1), .output_share0(d3_P1_13_s0), .output_share1(d3_P1_13_s1));
  reg_module u_reg_P1_17_d3 (.clk(clk), .input_share0(d2_P1_17_s0), .input_share1(d2_P1_17_s1), .output_share0(d3_P1_17_s0), .output_share1(d3_P1_17_s1));
  reg_module u_reg_P1_21_d3 (.clk(clk), .input_share0(d2_P1_21_s0), .input_share1(d2_P1_21_s1), .output_share0(d3_P1_21_s0), .output_share1(d3_P1_21_s1));
  reg_module u_reg_P1_25_d3 (.clk(clk), .input_share0(d2_P1_25_s0), .input_share1(d2_P1_25_s1), .output_share0(d3_P1_25_s0), .output_share1(d3_P1_25_s1));
  reg_module u_reg_P1_29_d3 (.clk(clk), .input_share0(d2_P1_29_s0), .input_share1(d2_P1_29_s1), .output_share0(d3_P1_29_s0), .output_share1(d3_P1_29_s1));
  reg_module u_reg_P1_5_d3 (.clk(clk), .input_share0(d2_P1_5_s0), .input_share1(d2_P1_5_s1), .output_share0(d3_P1_5_s0), .output_share1(d3_P1_5_s1));
  reg_module u_reg_P1_9_d3 (.clk(clk), .input_share0(d2_P1_9_s0), .input_share1(d2_P1_9_s1), .output_share0(d3_P1_9_s0), .output_share1(d3_P1_9_s1));
  reg_module u_reg_P2_10_d3 (.clk(clk), .input_share0(d2_P2_10_s0), .input_share1(d2_P2_10_s1), .output_share0(d3_P2_10_s0), .output_share1(d3_P2_10_s1));
  reg_module u_reg_P2_11_d3 (.clk(clk), .input_share0(d2_P2_11_s0), .input_share1(d2_P2_11_s1), .output_share0(d3_P2_11_s0), .output_share1(d3_P2_11_s1));
  reg_module u_reg_P2_14_d3 (.clk(clk), .input_share0(d2_P2_14_s0), .input_share1(d2_P2_14_s1), .output_share0(d3_P2_14_s0), .output_share1(d3_P2_14_s1));
  reg_module u_reg_P2_15_d3 (.clk(clk), .input_share0(d2_P2_15_s0), .input_share1(d2_P2_15_s1), .output_share0(d3_P2_15_s0), .output_share1(d3_P2_15_s1));
  reg_module u_reg_P2_18_d3 (.clk(clk), .input_share0(d2_P2_18_s0), .input_share1(d2_P2_18_s1), .output_share0(d3_P2_18_s0), .output_share1(d3_P2_18_s1));
  reg_module u_reg_P2_19_d3 (.clk(clk), .input_share0(d2_P2_19_s0), .input_share1(d2_P2_19_s1), .output_share0(d3_P2_19_s0), .output_share1(d3_P2_19_s1));
  reg_module u_reg_P2_22_d3 (.clk(clk), .input_share0(d2_P2_22_s0), .input_share1(d2_P2_22_s1), .output_share0(d3_P2_22_s0), .output_share1(d3_P2_22_s1));
  reg_module u_reg_P2_23_d3 (.clk(clk), .input_share0(d2_P2_23_s0), .input_share1(d2_P2_23_s1), .output_share0(d3_P2_23_s0), .output_share1(d3_P2_23_s1));
  reg_module u_reg_P2_26_d3 (.clk(clk), .input_share0(d2_P2_26_s0), .input_share1(d2_P2_26_s1), .output_share0(d3_P2_26_s0), .output_share1(d3_P2_26_s1));
  reg_module u_reg_P2_27_d3 (.clk(clk), .input_share0(d2_P2_27_s0), .input_share1(d2_P2_27_s1), .output_share0(d3_P2_27_s0), .output_share1(d3_P2_27_s1));
  reg_module u_reg_P2_30_d3 (.clk(clk), .input_share0(d2_P2_30_s0), .input_share1(d2_P2_30_s1), .output_share0(d3_P2_30_s0), .output_share1(d3_P2_30_s1));
  reg_module u_reg_P2_31_d3 (.clk(clk), .input_share0(d2_P2_31_s0), .input_share1(d2_P2_31_s1), .output_share0(d3_P2_31_s0), .output_share1(d3_P2_31_s1));
  reg_module u_reg_P2_6_d3 (.clk(clk), .input_share0(d2_P2_6_s0), .input_share1(d2_P2_6_s1), .output_share0(d3_P2_6_s0), .output_share1(d3_P2_6_s1));
  reg_module u_reg_P2_7_d3 (.clk(clk), .input_share0(d2_P2_7_s0), .input_share1(d2_P2_7_s1), .output_share0(d3_P2_7_s0), .output_share1(d3_P2_7_s1));
  xor_module u_xor_G2_10_d3 (.x_share0(d3_t20_s0), .x_share1(d3_t20_s1), .y_share0(d3_G0_10_s0), .y_share1(d3_G0_10_s1), .z_share0(d3_G2_10_s0), .z_share1(d3_G2_10_s1));
  xor_module u_xor_G2_11_d3 (.x_share0(d3_t21_s0), .x_share1(d3_t21_s1), .y_share0(d3_G1_11_s0), .y_share1(d3_G1_11_s1), .z_share0(d3_G2_11_s0), .z_share1(d3_G2_11_s1));
  xor_module u_xor_G2_14_d3 (.x_share0(d3_t22_s0), .x_share1(d3_t22_s1), .y_share0(d3_G0_14_s0), .y_share1(d3_G0_14_s1), .z_share0(d3_G2_14_s0), .z_share1(d3_G2_14_s1));
  xor_module u_xor_G2_15_d3 (.x_share0(d3_t23_s0), .x_share1(d3_t23_s1), .y_share0(d3_G1_15_s0), .y_share1(d3_G1_15_s1), .z_share0(d3_G2_15_s0), .z_share1(d3_G2_15_s1));
  xor_module u_xor_G2_18_d3 (.x_share0(d3_t24_s0), .x_share1(d3_t24_s1), .y_share0(d3_G0_18_s0), .y_share1(d3_G0_18_s1), .z_share0(d3_G2_18_s0), .z_share1(d3_G2_18_s1));
  xor_module u_xor_G2_19_d3 (.x_share0(d3_t25_s0), .x_share1(d3_t25_s1), .y_share0(d3_G1_19_s0), .y_share1(d3_G1_19_s1), .z_share0(d3_G2_19_s0), .z_share1(d3_G2_19_s1));
  xor_module u_xor_G2_2_d3 (.x_share0(d3_t16_s0), .x_share1(d3_t16_s1), .y_share0(d3_G0_2_s0), .y_share1(d3_G0_2_s1), .z_share0(d3_G2_2_s0), .z_share1(d3_G2_2_s1));
  xor_module u_xor_G2_22_d3 (.x_share0(d3_t26_s0), .x_share1(d3_t26_s1), .y_share0(d3_G0_22_s0), .y_share1(d3_G0_22_s1), .z_share0(d3_G2_22_s0), .z_share1(d3_G2_22_s1));
  xor_module u_xor_G2_23_d3 (.x_share0(d3_t27_s0), .x_share1(d3_t27_s1), .y_share0(d3_G1_23_s0), .y_share1(d3_G1_23_s1), .z_share0(d3_G2_23_s0), .z_share1(d3_G2_23_s1));
  xor_module u_xor_G2_26_d3 (.x_share0(d3_t28_s0), .x_share1(d3_t28_s1), .y_share0(d3_G0_26_s0), .y_share1(d3_G0_26_s1), .z_share0(d3_G2_26_s0), .z_share1(d3_G2_26_s1));
  xor_module u_xor_G2_27_d3 (.x_share0(d3_t29_s0), .x_share1(d3_t29_s1), .y_share0(d3_G1_27_s0), .y_share1(d3_G1_27_s1), .z_share0(d3_G2_27_s0), .z_share1(d3_G2_27_s1));
  xor_module u_xor_G2_3_d3 (.x_share0(d3_t17_s0), .x_share1(d3_t17_s1), .y_share0(d3_G1_3_s0), .y_share1(d3_G1_3_s1), .z_share0(d3_G2_3_s0), .z_share1(d3_G2_3_s1));
  xor_module u_xor_G2_30_d3 (.x_share0(d3_t30_s0), .x_share1(d3_t30_s1), .y_share0(d3_G0_30_s0), .y_share1(d3_G0_30_s1), .z_share0(d3_G2_30_s0), .z_share1(d3_G2_30_s1));
  xor_module u_xor_G2_31_d3 (.x_share0(d3_t31_s0), .x_share1(d3_t31_s1), .y_share0(d3_G1_31_s0), .y_share1(d3_G1_31_s1), .z_share0(d3_G2_31_s0), .z_share1(d3_G2_31_s1));
  xor_module u_xor_G2_6_d3 (.x_share0(d3_t18_s0), .x_share1(d3_t18_s1), .y_share0(d3_G0_6_s0), .y_share1(d3_G0_6_s1), .z_share0(d3_G2_6_s0), .z_share1(d3_G2_6_s1));
  xor_module u_xor_G2_7_d3 (.x_share0(d3_t19_s0), .x_share1(d3_t19_s1), .y_share0(d3_G1_7_s0), .y_share1(d3_G1_7_s1), .z_share0(d3_G2_7_s0), .z_share1(d3_G2_7_s1));
  and_module u_and_P3_12_d3 (.clk(clk), .x_share0(d2_P0_12_s0), .x_share1(d2_P0_12_s1), .y_share0(d2_P2_11_s0), .y_share1(d2_P2_11_s1), .rand(r_P3_12), .z_share0(d3_P3_12_s0), .z_share1(d3_P3_12_s1));
  assign r_P3_12 = stage3_share0[0];
  and_module u_and_P3_13_d3 (.clk(clk), .x_share0(d2_P1_13_s0), .x_share1(d2_P1_13_s1), .y_share0(d2_P2_11_s0), .y_share1(d2_P2_11_s1), .rand(r_P3_13), .z_share0(d3_P3_13_s0), .z_share1(d3_P3_13_s1));
  assign r_P3_13 = stage3_share0[2];
  and_module u_and_P3_14_d3 (.clk(clk), .x_share0(d2_P2_14_s0), .x_share1(d2_P2_14_s1), .y_share0(d2_P2_11_s0), .y_share1(d2_P2_11_s1), .rand(r_P3_14), .z_share0(d3_P3_14_s0), .z_share1(d3_P3_14_s1));
  assign r_P3_14 = stage3_share0[2];
  and_module u_and_P3_15_d3 (.clk(clk), .x_share0(d2_P2_15_s0), .x_share1(d2_P2_15_s1), .y_share0(d2_P2_11_s0), .y_share1(d2_P2_11_s1), .rand(r_P3_15), .z_share0(d3_P3_15_s0), .z_share1(d3_P3_15_s1));
  assign r_P3_15 = stage3_share0[2];
  and_module u_and_P3_20_d3 (.clk(clk), .x_share0(d2_P0_20_s0), .x_share1(d2_P0_20_s1), .y_share0(d2_P2_19_s0), .y_share1(d2_P2_19_s1), .rand(r_P3_20), .z_share0(d3_P3_20_s0), .z_share1(d3_P3_20_s1));
  assign r_P3_20 = stage3_share0[14];
  and_module u_and_P3_21_d3 (.clk(clk), .x_share0(d2_P1_21_s0), .x_share1(d2_P1_21_s1), .y_share0(d2_P2_19_s0), .y_share1(d2_P2_19_s1), .rand(r_P3_21), .z_share0(d3_P3_21_s0), .z_share1(d3_P3_21_s1));
  assign r_P3_21 = stage3_share0[14];
  and_module u_and_P3_22_d3 (.clk(clk), .x_share0(d2_P2_22_s0), .x_share1(d2_P2_22_s1), .y_share0(d2_P2_19_s0), .y_share1(d2_P2_19_s1), .rand(r_P3_22), .z_share0(d3_P3_22_s0), .z_share1(d3_P3_22_s1));
  assign r_P3_22 = stage3_share0[15];
  and_module u_and_P3_23_d3 (.clk(clk), .x_share0(d2_P2_23_s0), .x_share1(d2_P2_23_s1), .y_share0(d2_P2_19_s0), .y_share1(d2_P2_19_s1), .rand(r_P3_23), .z_share0(d3_P3_23_s0), .z_share1(d3_P3_23_s1));
  assign r_P3_23 = stage3_share0[22];
  and_module u_and_P3_28_d3 (.clk(clk), .x_share0(d2_P0_28_s0), .x_share1(d2_P0_28_s1), .y_share0(d2_P2_27_s0), .y_share1(d2_P2_27_s1), .rand(r_P3_28), .z_share0(d3_P3_28_s0), .z_share1(d3_P3_28_s1));
  assign r_P3_28 = stage3_share0[19];
  and_module u_and_P3_29_d3 (.clk(clk), .x_share0(d2_P1_29_s0), .x_share1(d2_P1_29_s1), .y_share0(d2_P2_27_s0), .y_share1(d2_P2_27_s1), .rand(r_P3_29), .z_share0(d3_P3_29_s0), .z_share1(d3_P3_29_s1));
  assign r_P3_29 = stage3_share0[19];
  and_module u_and_P3_30_d3 (.clk(clk), .x_share0(d2_P2_30_s0), .x_share1(d2_P2_30_s1), .y_share0(d2_P2_27_s0), .y_share1(d2_P2_27_s1), .rand(r_P3_30), .z_share0(d3_P3_30_s0), .z_share1(d3_P3_30_s1));
  assign r_P3_30 = stage3_share0[23];
  and_module u_and_P3_31_d3 (.clk(clk), .x_share0(d2_P2_31_s0), .x_share1(d2_P2_31_s1), .y_share0(d2_P2_27_s0), .y_share1(d2_P2_27_s1), .rand(r_P3_31), .z_share0(d3_P3_31_s0), .z_share1(d3_P3_31_s1));
  assign r_P3_31 = stage3_share0[25];
  xor_module u_xor_o3_d3 (.x_share0(d3_P0_3_s0), .x_share1(d3_P0_3_s1), .y_share0(d3_G2_2_s0), .y_share1(d3_G2_2_s1), .z_share0(d3_o3_s0), .z_share1(d3_o3_s1));
  xor_module u_xor_o4_d3 (.x_share0(d3_P0_4_s0), .x_share1(d3_P0_4_s1), .y_share0(d3_G2_3_s0), .y_share1(d3_G2_3_s1), .z_share0(d3_o4_s0), .z_share1(d3_o4_s1));
  and_module u_and_t16_d3 (.clk(clk), .x_share0(d2_P0_2_s0), .x_share1(d2_P0_2_s1), .y_share0(d2_G1_1_s0), .y_share1(d2_G1_1_s1), .rand(r_t16), .z_share0(d3_t16_s0), .z_share1(d3_t16_s1));
  assign r_t16 = stage3_share0[3];
  and_module u_and_t17_d3 (.clk(clk), .x_share0(d2_P1_3_s0), .x_share1(d2_P1_3_s1), .y_share0(d2_G1_1_s0), .y_share1(d2_G1_1_s1), .rand(r_t17), .z_share0(d3_t17_s0), .z_share1(d3_t17_s1));
  assign r_t17 = stage3_share0[16];
  and_module u_and_t18_d3 (.clk(clk), .x_share0(d2_P0_6_s0), .x_share1(d2_P0_6_s1), .y_share0(d2_G1_5_s0), .y_share1(d2_G1_5_s1), .rand(r_t18), .z_share0(d3_t18_s0), .z_share1(d3_t18_s1));
  assign r_t18 = stage3_share0[4];
  and_module u_and_t19_d3 (.clk(clk), .x_share0(d2_P1_7_s0), .x_share1(d2_P1_7_s1), .y_share0(d2_G1_5_s0), .y_share1(d2_G1_5_s1), .rand(r_t19), .z_share0(d3_t19_s0), .z_share1(d3_t19_s1));
  assign r_t19 = stage3_share0[12];
  and_module u_and_t20_d3 (.clk(clk), .x_share0(d2_P0_10_s0), .x_share1(d2_P0_10_s1), .y_share0(d2_G1_9_s0), .y_share1(d2_G1_9_s1), .rand(r_t20), .z_share0(d3_t20_s0), .z_share1(d3_t20_s1));
  assign r_t20 = stage3_share0[3];
  and_module u_and_t21_d3 (.clk(clk), .x_share0(d2_P1_11_s0), .x_share1(d2_P1_11_s1), .y_share0(d2_G1_9_s0), .y_share1(d2_G1_9_s1), .rand(r_t21), .z_share0(d3_t21_s0), .z_share1(d3_t21_s1));
  assign r_t21 = stage3_share0[15];
  and_module u_and_t22_d3 (.clk(clk), .x_share0(d2_P0_14_s0), .x_share1(d2_P0_14_s1), .y_share0(d2_G1_13_s0), .y_share1(d2_G1_13_s1), .rand(r_t22), .z_share0(d3_t22_s0), .z_share1(d3_t22_s1));
  assign r_t22 = stage3_share0[4];
  and_module u_and_t23_d3 (.clk(clk), .x_share0(d2_P1_15_s0), .x_share1(d2_P1_15_s1), .y_share0(d2_G1_13_s0), .y_share1(d2_G1_13_s1), .rand(r_t23), .z_share0(d3_t23_s0), .z_share1(d3_t23_s1));
  assign r_t23 = stage3_share0[5];
  and_module u_and_t24_d3 (.clk(clk), .x_share0(d2_P0_18_s0), .x_share1(d2_P0_18_s1), .y_share0(d2_G1_17_s0), .y_share1(d2_G1_17_s1), .rand(r_t24), .z_share0(d3_t24_s0), .z_share1(d3_t24_s1));
  assign r_t24 = stage3_share0[11];
  and_module u_and_t25_d3 (.clk(clk), .x_share0(d2_P1_19_s0), .x_share1(d2_P1_19_s1), .y_share0(d2_G1_17_s0), .y_share1(d2_G1_17_s1), .rand(r_t25), .z_share0(d3_t25_s0), .z_share1(d3_t25_s1));
  assign r_t25 = stage3_share0[22];
  and_module u_and_t26_d3 (.clk(clk), .x_share0(d2_P0_22_s0), .x_share1(d2_P0_22_s1), .y_share0(d2_G1_21_s0), .y_share1(d2_G1_21_s1), .rand(r_t26), .z_share0(d3_t26_s0), .z_share1(d3_t26_s1));
  assign r_t26 = stage3_share0[9];
  and_module u_and_t27_d3 (.clk(clk), .x_share0(d2_P1_23_s0), .x_share1(d2_P1_23_s1), .y_share0(d2_G1_21_s0), .y_share1(d2_G1_21_s1), .rand(r_t27), .z_share0(d3_t27_s0), .z_share1(d3_t27_s1));
  assign r_t27 = stage3_share0[10];
  and_module u_and_t28_d3 (.clk(clk), .x_share0(d2_P0_26_s0), .x_share1(d2_P0_26_s1), .y_share0(d2_G1_25_s0), .y_share1(d2_G1_25_s1), .rand(r_t28), .z_share0(d3_t28_s0), .z_share1(d3_t28_s1));
  assign r_t28 = stage3_share0[12];
  and_module u_and_t29_d3 (.clk(clk), .x_share0(d2_P1_27_s0), .x_share1(d2_P1_27_s1), .y_share0(d2_G1_25_s0), .y_share1(d2_G1_25_s1), .rand(r_t29), .z_share0(d3_t29_s0), .z_share1(d3_t29_s1));
  assign r_t29 = stage3_share0[16];
  and_module u_and_t30_d3 (.clk(clk), .x_share0(d2_P0_30_s0), .x_share1(d2_P0_30_s1), .y_share0(d2_G1_29_s0), .y_share1(d2_G1_29_s1), .rand(r_t30), .z_share0(d3_t30_s0), .z_share1(d3_t30_s1));
  assign r_t30 = stage3_share0[18];
  and_module u_and_t31_d3 (.clk(clk), .x_share0(d2_P1_31_s0), .x_share1(d2_P1_31_s1), .y_share0(d2_G1_29_s0), .y_share1(d2_G1_29_s1), .rand(r_t31), .z_share0(d3_t31_s0), .z_share1(d3_t31_s1));
  assign r_t31 = stage3_share0[24];
  reg_module u_reg_G0_12_d4 (.clk(clk), .input_share0(d3_G0_12_s0), .input_share1(d3_G0_12_s1), .output_share0(d4_G0_12_s0), .output_share1(d4_G0_12_s1));
  reg_module u_reg_G0_16_d4 (.clk(clk), .input_share0(d3_G0_16_s0), .input_share1(d3_G0_16_s1), .output_share0(d4_G0_16_s0), .output_share1(d4_G0_16_s1));
  reg_module u_reg_G0_20_d4 (.clk(clk), .input_share0(d3_G0_20_s0), .input_share1(d3_G0_20_s1), .output_share0(d4_G0_20_s0), .output_share1(d4_G0_20_s1));
  reg_module u_reg_G0_24_d4 (.clk(clk), .input_share0(d3_G0_24_s0), .input_share1(d3_G0_24_s1), .output_share0(d4_G0_24_s0), .output_share1(d4_G0_24_s1));
  reg_module u_reg_G0_28_d4 (.clk(clk), .input_share0(d3_G0_28_s0), .input_share1(d3_G0_28_s1), .output_share0(d4_G0_28_s0), .output_share1(d4_G0_28_s1));
  reg_module u_reg_G0_4_d4 (.clk(clk), .input_share0(d3_G0_4_s0), .input_share1(d3_G0_4_s1), .output_share0(d4_G0_4_s0), .output_share1(d4_G0_4_s1));
  reg_module u_reg_G0_8_d4 (.clk(clk), .input_share0(d3_G0_8_s0), .input_share1(d3_G0_8_s1), .output_share0(d4_G0_8_s0), .output_share1(d4_G0_8_s1));
  reg_module u_reg_G1_13_d4 (.clk(clk), .input_share0(d3_G1_13_s0), .input_share1(d3_G1_13_s1), .output_share0(d4_G1_13_s0), .output_share1(d4_G1_13_s1));
  reg_module u_reg_G1_17_d4 (.clk(clk), .input_share0(d3_G1_17_s0), .input_share1(d3_G1_17_s1), .output_share0(d4_G1_17_s0), .output_share1(d4_G1_17_s1));
  reg_module u_reg_G1_21_d4 (.clk(clk), .input_share0(d3_G1_21_s0), .input_share1(d3_G1_21_s1), .output_share0(d4_G1_21_s0), .output_share1(d4_G1_21_s1));
  reg_module u_reg_G1_25_d4 (.clk(clk), .input_share0(d3_G1_25_s0), .input_share1(d3_G1_25_s1), .output_share0(d4_G1_25_s0), .output_share1(d4_G1_25_s1));
  reg_module u_reg_G1_29_d4 (.clk(clk), .input_share0(d3_G1_29_s0), .input_share1(d3_G1_29_s1), .output_share0(d4_G1_29_s0), .output_share1(d4_G1_29_s1));
  reg_module u_reg_G1_5_d4 (.clk(clk), .input_share0(d3_G1_5_s0), .input_share1(d3_G1_5_s1), .output_share0(d4_G1_5_s0), .output_share1(d4_G1_5_s1));
  reg_module u_reg_G1_9_d4 (.clk(clk), .input_share0(d3_G1_9_s0), .input_share1(d3_G1_9_s1), .output_share0(d4_G1_9_s0), .output_share1(d4_G1_9_s1));
  reg_module u_reg_G2_10_d4 (.clk(clk), .input_share0(d3_G2_10_s0), .input_share1(d3_G2_10_s1), .output_share0(d4_G2_10_s0), .output_share1(d4_G2_10_s1));
  reg_module u_reg_G2_11_d4 (.clk(clk), .input_share0(d3_G2_11_s0), .input_share1(d3_G2_11_s1), .output_share0(d4_G2_11_s0), .output_share1(d4_G2_11_s1));
  reg_module u_reg_G2_14_d4 (.clk(clk), .input_share0(d3_G2_14_s0), .input_share1(d3_G2_14_s1), .output_share0(d4_G2_14_s0), .output_share1(d4_G2_14_s1));
  reg_module u_reg_G2_15_d4 (.clk(clk), .input_share0(d3_G2_15_s0), .input_share1(d3_G2_15_s1), .output_share0(d4_G2_15_s0), .output_share1(d4_G2_15_s1));
  reg_module u_reg_G2_18_d4 (.clk(clk), .input_share0(d3_G2_18_s0), .input_share1(d3_G2_18_s1), .output_share0(d4_G2_18_s0), .output_share1(d4_G2_18_s1));
  reg_module u_reg_G2_19_d4 (.clk(clk), .input_share0(d3_G2_19_s0), .input_share1(d3_G2_19_s1), .output_share0(d4_G2_19_s0), .output_share1(d4_G2_19_s1));
  reg_module u_reg_G2_22_d4 (.clk(clk), .input_share0(d3_G2_22_s0), .input_share1(d3_G2_22_s1), .output_share0(d4_G2_22_s0), .output_share1(d4_G2_22_s1));
  reg_module u_reg_G2_23_d4 (.clk(clk), .input_share0(d3_G2_23_s0), .input_share1(d3_G2_23_s1), .output_share0(d4_G2_23_s0), .output_share1(d4_G2_23_s1));
  reg_module u_reg_G2_26_d4 (.clk(clk), .input_share0(d3_G2_26_s0), .input_share1(d3_G2_26_s1), .output_share0(d4_G2_26_s0), .output_share1(d4_G2_26_s1));
  reg_module u_reg_G2_27_d4 (.clk(clk), .input_share0(d3_G2_27_s0), .input_share1(d3_G2_27_s1), .output_share0(d4_G2_27_s0), .output_share1(d4_G2_27_s1));
  reg_module u_reg_G2_30_d4 (.clk(clk), .input_share0(d3_G2_30_s0), .input_share1(d3_G2_30_s1), .output_share0(d4_G2_30_s0), .output_share1(d4_G2_30_s1));
  reg_module u_reg_G2_31_d4 (.clk(clk), .input_share0(d3_G2_31_s0), .input_share1(d3_G2_31_s1), .output_share0(d4_G2_31_s0), .output_share1(d4_G2_31_s1));
  reg_module u_reg_G2_6_d4 (.clk(clk), .input_share0(d3_G2_6_s0), .input_share1(d3_G2_6_s1), .output_share0(d4_G2_6_s0), .output_share1(d4_G2_6_s1));
  reg_module u_reg_G2_7_d4 (.clk(clk), .input_share0(d3_G2_7_s0), .input_share1(d3_G2_7_s1), .output_share0(d4_G2_7_s0), .output_share1(d4_G2_7_s1));
  reg_module u_reg_P0_10_d4 (.clk(clk), .input_share0(d3_P0_10_s0), .input_share1(d3_P0_10_s1), .output_share0(d4_P0_10_s0), .output_share1(d4_P0_10_s1));
  reg_module u_reg_P0_11_d4 (.clk(clk), .input_share0(d3_P0_11_s0), .input_share1(d3_P0_11_s1), .output_share0(d4_P0_11_s0), .output_share1(d4_P0_11_s1));
  reg_module u_reg_P0_12_d4 (.clk(clk), .input_share0(d3_P0_12_s0), .input_share1(d3_P0_12_s1), .output_share0(d4_P0_12_s0), .output_share1(d4_P0_12_s1));
  reg_module u_reg_P0_13_d4 (.clk(clk), .input_share0(d3_P0_13_s0), .input_share1(d3_P0_13_s1), .output_share0(d4_P0_13_s0), .output_share1(d4_P0_13_s1));
  reg_module u_reg_P0_14_d4 (.clk(clk), .input_share0(d3_P0_14_s0), .input_share1(d3_P0_14_s1), .output_share0(d4_P0_14_s0), .output_share1(d4_P0_14_s1));
  reg_module u_reg_P0_15_d4 (.clk(clk), .input_share0(d3_P0_15_s0), .input_share1(d3_P0_15_s1), .output_share0(d4_P0_15_s0), .output_share1(d4_P0_15_s1));
  reg_module u_reg_P0_16_d4 (.clk(clk), .input_share0(d3_P0_16_s0), .input_share1(d3_P0_16_s1), .output_share0(d4_P0_16_s0), .output_share1(d4_P0_16_s1));
  reg_module u_reg_P0_17_d4 (.clk(clk), .input_share0(d3_P0_17_s0), .input_share1(d3_P0_17_s1), .output_share0(d4_P0_17_s0), .output_share1(d4_P0_17_s1));
  reg_module u_reg_P0_18_d4 (.clk(clk), .input_share0(d3_P0_18_s0), .input_share1(d3_P0_18_s1), .output_share0(d4_P0_18_s0), .output_share1(d4_P0_18_s1));
  reg_module u_reg_P0_19_d4 (.clk(clk), .input_share0(d3_P0_19_s0), .input_share1(d3_P0_19_s1), .output_share0(d4_P0_19_s0), .output_share1(d4_P0_19_s1));
  reg_module u_reg_P0_20_d4 (.clk(clk), .input_share0(d3_P0_20_s0), .input_share1(d3_P0_20_s1), .output_share0(d4_P0_20_s0), .output_share1(d4_P0_20_s1));
  reg_module u_reg_P0_21_d4 (.clk(clk), .input_share0(d3_P0_21_s0), .input_share1(d3_P0_21_s1), .output_share0(d4_P0_21_s0), .output_share1(d4_P0_21_s1));
  reg_module u_reg_P0_22_d4 (.clk(clk), .input_share0(d3_P0_22_s0), .input_share1(d3_P0_22_s1), .output_share0(d4_P0_22_s0), .output_share1(d4_P0_22_s1));
  reg_module u_reg_P0_23_d4 (.clk(clk), .input_share0(d3_P0_23_s0), .input_share1(d3_P0_23_s1), .output_share0(d4_P0_23_s0), .output_share1(d4_P0_23_s1));
  reg_module u_reg_P0_24_d4 (.clk(clk), .input_share0(d3_P0_24_s0), .input_share1(d3_P0_24_s1), .output_share0(d4_P0_24_s0), .output_share1(d4_P0_24_s1));
  reg_module u_reg_P0_25_d4 (.clk(clk), .input_share0(d3_P0_25_s0), .input_share1(d3_P0_25_s1), .output_share0(d4_P0_25_s0), .output_share1(d4_P0_25_s1));
  reg_module u_reg_P0_26_d4 (.clk(clk), .input_share0(d3_P0_26_s0), .input_share1(d3_P0_26_s1), .output_share0(d4_P0_26_s0), .output_share1(d4_P0_26_s1));
  reg_module u_reg_P0_27_d4 (.clk(clk), .input_share0(d3_P0_27_s0), .input_share1(d3_P0_27_s1), .output_share0(d4_P0_27_s0), .output_share1(d4_P0_27_s1));
  reg_module u_reg_P0_28_d4 (.clk(clk), .input_share0(d3_P0_28_s0), .input_share1(d3_P0_28_s1), .output_share0(d4_P0_28_s0), .output_share1(d4_P0_28_s1));
  reg_module u_reg_P0_29_d4 (.clk(clk), .input_share0(d3_P0_29_s0), .input_share1(d3_P0_29_s1), .output_share0(d4_P0_29_s0), .output_share1(d4_P0_29_s1));
  reg_module u_reg_P0_30_d4 (.clk(clk), .input_share0(d3_P0_30_s0), .input_share1(d3_P0_30_s1), .output_share0(d4_P0_30_s0), .output_share1(d4_P0_30_s1));
  reg_module u_reg_P0_31_d4 (.clk(clk), .input_share0(d3_P0_31_s0), .input_share1(d3_P0_31_s1), .output_share0(d4_P0_31_s0), .output_share1(d4_P0_31_s1));
  reg_module u_reg_P0_5_d4 (.clk(clk), .input_share0(d3_P0_5_s0), .input_share1(d3_P0_5_s1), .output_share0(d4_P0_5_s0), .output_share1(d4_P0_5_s1));
  reg_module u_reg_P0_6_d4 (.clk(clk), .input_share0(d3_P0_6_s0), .input_share1(d3_P0_6_s1), .output_share0(d4_P0_6_s0), .output_share1(d4_P0_6_s1));
  reg_module u_reg_P0_7_d4 (.clk(clk), .input_share0(d3_P0_7_s0), .input_share1(d3_P0_7_s1), .output_share0(d4_P0_7_s0), .output_share1(d4_P0_7_s1));
  reg_module u_reg_P0_8_d4 (.clk(clk), .input_share0(d3_P0_8_s0), .input_share1(d3_P0_8_s1), .output_share0(d4_P0_8_s0), .output_share1(d4_P0_8_s1));
  reg_module u_reg_P0_9_d4 (.clk(clk), .input_share0(d3_P0_9_s0), .input_share1(d3_P0_9_s1), .output_share0(d4_P0_9_s0), .output_share1(d4_P0_9_s1));
  reg_module u_reg_P1_17_d4 (.clk(clk), .input_share0(d3_P1_17_s0), .input_share1(d3_P1_17_s1), .output_share0(d4_P1_17_s0), .output_share1(d4_P1_17_s1));
  reg_module u_reg_P1_25_d4 (.clk(clk), .input_share0(d3_P1_25_s0), .input_share1(d3_P1_25_s1), .output_share0(d4_P1_25_s0), .output_share1(d4_P1_25_s1));
  reg_module u_reg_P1_9_d4 (.clk(clk), .input_share0(d3_P1_9_s0), .input_share1(d3_P1_9_s1), .output_share0(d4_P1_9_s0), .output_share1(d4_P1_9_s1));
  reg_module u_reg_P2_10_d4 (.clk(clk), .input_share0(d3_P2_10_s0), .input_share1(d3_P2_10_s1), .output_share0(d4_P2_10_s0), .output_share1(d4_P2_10_s1));
  reg_module u_reg_P2_11_d4 (.clk(clk), .input_share0(d3_P2_11_s0), .input_share1(d3_P2_11_s1), .output_share0(d4_P2_11_s0), .output_share1(d4_P2_11_s1));
  reg_module u_reg_P2_18_d4 (.clk(clk), .input_share0(d3_P2_18_s0), .input_share1(d3_P2_18_s1), .output_share0(d4_P2_18_s0), .output_share1(d4_P2_18_s1));
  reg_module u_reg_P2_19_d4 (.clk(clk), .input_share0(d3_P2_19_s0), .input_share1(d3_P2_19_s1), .output_share0(d4_P2_19_s0), .output_share1(d4_P2_19_s1));
  reg_module u_reg_P2_26_d4 (.clk(clk), .input_share0(d3_P2_26_s0), .input_share1(d3_P2_26_s1), .output_share0(d4_P2_26_s0), .output_share1(d4_P2_26_s1));
  reg_module u_reg_P2_27_d4 (.clk(clk), .input_share0(d3_P2_27_s0), .input_share1(d3_P2_27_s1), .output_share0(d4_P2_27_s0), .output_share1(d4_P2_27_s1));
  reg_module u_reg_P3_12_d4 (.clk(clk), .input_share0(d3_P3_12_s0), .input_share1(d3_P3_12_s1), .output_share0(d4_P3_12_s0), .output_share1(d4_P3_12_s1));
  reg_module u_reg_P3_13_d4 (.clk(clk), .input_share0(d3_P3_13_s0), .input_share1(d3_P3_13_s1), .output_share0(d4_P3_13_s0), .output_share1(d4_P3_13_s1));
  reg_module u_reg_P3_14_d4 (.clk(clk), .input_share0(d3_P3_14_s0), .input_share1(d3_P3_14_s1), .output_share0(d4_P3_14_s0), .output_share1(d4_P3_14_s1));
  reg_module u_reg_P3_15_d4 (.clk(clk), .input_share0(d3_P3_15_s0), .input_share1(d3_P3_15_s1), .output_share0(d4_P3_15_s0), .output_share1(d4_P3_15_s1));
  reg_module u_reg_P3_20_d4 (.clk(clk), .input_share0(d3_P3_20_s0), .input_share1(d3_P3_20_s1), .output_share0(d4_P3_20_s0), .output_share1(d4_P3_20_s1));
  reg_module u_reg_P3_21_d4 (.clk(clk), .input_share0(d3_P3_21_s0), .input_share1(d3_P3_21_s1), .output_share0(d4_P3_21_s0), .output_share1(d4_P3_21_s1));
  reg_module u_reg_P3_22_d4 (.clk(clk), .input_share0(d3_P3_22_s0), .input_share1(d3_P3_22_s1), .output_share0(d4_P3_22_s0), .output_share1(d4_P3_22_s1));
  reg_module u_reg_P3_23_d4 (.clk(clk), .input_share0(d3_P3_23_s0), .input_share1(d3_P3_23_s1), .output_share0(d4_P3_23_s0), .output_share1(d4_P3_23_s1));
  reg_module u_reg_P3_28_d4 (.clk(clk), .input_share0(d3_P3_28_s0), .input_share1(d3_P3_28_s1), .output_share0(d4_P3_28_s0), .output_share1(d4_P3_28_s1));
  reg_module u_reg_P3_29_d4 (.clk(clk), .input_share0(d3_P3_29_s0), .input_share1(d3_P3_29_s1), .output_share0(d4_P3_29_s0), .output_share1(d4_P3_29_s1));
  reg_module u_reg_P3_30_d4 (.clk(clk), .input_share0(d3_P3_30_s0), .input_share1(d3_P3_30_s1), .output_share0(d4_P3_30_s0), .output_share1(d4_P3_30_s1));
  reg_module u_reg_P3_31_d4 (.clk(clk), .input_share0(d3_P3_31_s0), .input_share1(d3_P3_31_s1), .output_share0(d4_P3_31_s0), .output_share1(d4_P3_31_s1));
  xor_module u_xor_G3_12_d4 (.x_share0(d4_t36_s0), .x_share1(d4_t36_s1), .y_share0(d4_G0_12_s0), .y_share1(d4_G0_12_s1), .z_share0(d4_G3_12_s0), .z_share1(d4_G3_12_s1));
  xor_module u_xor_G3_13_d4 (.x_share0(d4_t37_s0), .x_share1(d4_t37_s1), .y_share0(d4_G1_13_s0), .y_share1(d4_G1_13_s1), .z_share0(d4_G3_13_s0), .z_share1(d4_G3_13_s1));
  xor_module u_xor_G3_14_d4 (.x_share0(d4_t38_s0), .x_share1(d4_t38_s1), .y_share0(d4_G2_14_s0), .y_share1(d4_G2_14_s1), .z_share0(d4_G3_14_s0), .z_share1(d4_G3_14_s1));
  xor_module u_xor_G3_15_d4 (.x_share0(d4_t39_s0), .x_share1(d4_t39_s1), .y_share0(d4_G2_15_s0), .y_share1(d4_G2_15_s1), .z_share0(d4_G3_15_s0), .z_share1(d4_G3_15_s1));
  xor_module u_xor_G3_20_d4 (.x_share0(d4_t40_s0), .x_share1(d4_t40_s1), .y_share0(d4_G0_20_s0), .y_share1(d4_G0_20_s1), .z_share0(d4_G3_20_s0), .z_share1(d4_G3_20_s1));
  xor_module u_xor_G3_21_d4 (.x_share0(d4_t41_s0), .x_share1(d4_t41_s1), .y_share0(d4_G1_21_s0), .y_share1(d4_G1_21_s1), .z_share0(d4_G3_21_s0), .z_share1(d4_G3_21_s1));
  xor_module u_xor_G3_22_d4 (.x_share0(d4_t42_s0), .x_share1(d4_t42_s1), .y_share0(d4_G2_22_s0), .y_share1(d4_G2_22_s1), .z_share0(d4_G3_22_s0), .z_share1(d4_G3_22_s1));
  xor_module u_xor_G3_23_d4 (.x_share0(d4_t43_s0), .x_share1(d4_t43_s1), .y_share0(d4_G2_23_s0), .y_share1(d4_G2_23_s1), .z_share0(d4_G3_23_s0), .z_share1(d4_G3_23_s1));
  xor_module u_xor_G3_28_d4 (.x_share0(d4_t44_s0), .x_share1(d4_t44_s1), .y_share0(d4_G0_28_s0), .y_share1(d4_G0_28_s1), .z_share0(d4_G3_28_s0), .z_share1(d4_G3_28_s1));
  xor_module u_xor_G3_29_d4 (.x_share0(d4_t45_s0), .x_share1(d4_t45_s1), .y_share0(d4_G1_29_s0), .y_share1(d4_G1_29_s1), .z_share0(d4_G3_29_s0), .z_share1(d4_G3_29_s1));
  xor_module u_xor_G3_30_d4 (.x_share0(d4_t46_s0), .x_share1(d4_t46_s1), .y_share0(d4_G2_30_s0), .y_share1(d4_G2_30_s1), .z_share0(d4_G3_30_s0), .z_share1(d4_G3_30_s1));
  xor_module u_xor_G3_31_d4 (.x_share0(d4_t47_s0), .x_share1(d4_t47_s1), .y_share0(d4_G2_31_s0), .y_share1(d4_G2_31_s1), .z_share0(d4_G3_31_s0), .z_share1(d4_G3_31_s1));
  xor_module u_xor_G3_4_d4 (.x_share0(d4_t32_s0), .x_share1(d4_t32_s1), .y_share0(d4_G0_4_s0), .y_share1(d4_G0_4_s1), .z_share0(d4_G3_4_s0), .z_share1(d4_G3_4_s1));
  xor_module u_xor_G3_5_d4 (.x_share0(d4_t33_s0), .x_share1(d4_t33_s1), .y_share0(d4_G1_5_s0), .y_share1(d4_G1_5_s1), .z_share0(d4_G3_5_s0), .z_share1(d4_G3_5_s1));
  xor_module u_xor_G3_6_d4 (.x_share0(d4_t34_s0), .x_share1(d4_t34_s1), .y_share0(d4_G2_6_s0), .y_share1(d4_G2_6_s1), .z_share0(d4_G3_6_s0), .z_share1(d4_G3_6_s1));
  xor_module u_xor_G3_7_d4 (.x_share0(d4_t35_s0), .x_share1(d4_t35_s1), .y_share0(d4_G2_7_s0), .y_share1(d4_G2_7_s1), .z_share0(d4_G3_7_s0), .z_share1(d4_G3_7_s1));
  and_module u_and_P4_24_d4 (.clk(clk), .x_share0(d3_P0_24_s0), .x_share1(d3_P0_24_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_24), .z_share0(d4_P4_24_s0), .z_share1(d4_P4_24_s1));
  assign r_P4_24 = stage4_share0[17];
  and_module u_and_P4_25_d4 (.clk(clk), .x_share0(d3_P1_25_s0), .x_share1(d3_P1_25_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_25), .z_share0(d4_P4_25_s0), .z_share1(d4_P4_25_s1));
  assign r_P4_25 = stage4_share0[17];
  and_module u_and_P4_26_d4 (.clk(clk), .x_share0(d3_P2_26_s0), .x_share1(d3_P2_26_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_26), .z_share0(d4_P4_26_s0), .z_share1(d4_P4_26_s1));
  assign r_P4_26 = stage4_share0[19];
  and_module u_and_P4_27_d4 (.clk(clk), .x_share0(d3_P2_27_s0), .x_share1(d3_P2_27_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_27), .z_share0(d4_P4_27_s0), .z_share1(d4_P4_27_s1));
  assign r_P4_27 = stage4_share0[19];
  and_module u_and_P4_28_d4 (.clk(clk), .x_share0(d3_P3_28_s0), .x_share1(d3_P3_28_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_28), .z_share0(d4_P4_28_s0), .z_share1(d4_P4_28_s1));
  assign r_P4_28 = stage4_share0[20];
  and_module u_and_P4_29_d4 (.clk(clk), .x_share0(d3_P3_29_s0), .x_share1(d3_P3_29_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_29), .z_share0(d4_P4_29_s0), .z_share1(d4_P4_29_s1));
  assign r_P4_29 = stage4_share0[23];
  and_module u_and_P4_30_d4 (.clk(clk), .x_share0(d3_P3_30_s0), .x_share1(d3_P3_30_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_30), .z_share0(d4_P4_30_s0), .z_share1(d4_P4_30_s1));
  assign r_P4_30 = stage4_share0[20];
  and_module u_and_P4_31_d4 (.clk(clk), .x_share0(d3_P3_31_s0), .x_share1(d3_P3_31_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_31), .z_share0(d4_P4_31_s0), .z_share1(d4_P4_31_s1));
  assign r_P4_31 = stage4_share0[20];
  xor_module u_xor_o5_d4 (.x_share0(d4_P0_5_s0), .x_share1(d4_P0_5_s1), .y_share0(d4_G3_4_s0), .y_share1(d4_G3_4_s1), .z_share0(d4_o5_s0), .z_share1(d4_o5_s1));
  xor_module u_xor_o6_d4 (.x_share0(d4_P0_6_s0), .x_share1(d4_P0_6_s1), .y_share0(d4_G3_5_s0), .y_share1(d4_G3_5_s1), .z_share0(d4_o6_s0), .z_share1(d4_o6_s1));
  xor_module u_xor_o7_d4 (.x_share0(d4_P0_7_s0), .x_share1(d4_P0_7_s1), .y_share0(d4_G3_6_s0), .y_share1(d4_G3_6_s1), .z_share0(d4_o7_s0), .z_share1(d4_o7_s1));
  xor_module u_xor_o8_d4 (.x_share0(d4_P0_8_s0), .x_share1(d4_P0_8_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .z_share0(d4_o8_s0), .z_share1(d4_o8_s1));
  and_module u_and_t32_d4 (.clk(clk), .x_share0(d3_P0_4_s0), .x_share1(d3_P0_4_s1), .y_share0(d3_G2_3_s0), .y_share1(d3_G2_3_s1), .rand(r_t32), .z_share0(d4_t32_s0), .z_share1(d4_t32_s1));
  assign r_t32 = stage4_share0[3];
  and_module u_and_t33_d4 (.clk(clk), .x_share0(d3_P1_5_s0), .x_share1(d3_P1_5_s1), .y_share0(d3_G2_3_s0), .y_share1(d3_G2_3_s1), .rand(r_t33), .z_share0(d4_t33_s0), .z_share1(d4_t33_s1));
  assign r_t33 = stage4_share0[3];
  and_module u_and_t34_d4 (.clk(clk), .x_share0(d3_P2_6_s0), .x_share1(d3_P2_6_s1), .y_share0(d3_G2_3_s0), .y_share1(d3_G2_3_s1), .rand(r_t34), .z_share0(d4_t34_s0), .z_share1(d4_t34_s1));
  assign r_t34 = stage4_share0[6];
  and_module u_and_t35_d4 (.clk(clk), .x_share0(d3_P2_7_s0), .x_share1(d3_P2_7_s1), .y_share0(d3_G2_3_s0), .y_share1(d3_G2_3_s1), .rand(r_t35), .z_share0(d4_t35_s0), .z_share1(d4_t35_s1));
  assign r_t35 = stage4_share0[13];
  and_module u_and_t36_d4 (.clk(clk), .x_share0(d3_P0_12_s0), .x_share1(d3_P0_12_s1), .y_share0(d3_G2_11_s0), .y_share1(d3_G2_11_s1), .rand(r_t36), .z_share0(d4_t36_s0), .z_share1(d4_t36_s1));
  assign r_t36 = stage4_share0[1];
  and_module u_and_t37_d4 (.clk(clk), .x_share0(d3_P1_13_s0), .x_share1(d3_P1_13_s1), .y_share0(d3_G2_11_s0), .y_share1(d3_G2_11_s1), .rand(r_t37), .z_share0(d4_t37_s0), .z_share1(d4_t37_s1));
  assign r_t37 = stage4_share0[0];
  and_module u_and_t38_d4 (.clk(clk), .x_share0(d3_P2_14_s0), .x_share1(d3_P2_14_s1), .y_share0(d3_G2_11_s0), .y_share1(d3_G2_11_s1), .rand(r_t38), .z_share0(d4_t38_s0), .z_share1(d4_t38_s1));
  assign r_t38 = stage4_share0[3];
  and_module u_and_t39_d4 (.clk(clk), .x_share0(d3_P2_15_s0), .x_share1(d3_P2_15_s1), .y_share0(d3_G2_11_s0), .y_share1(d3_G2_11_s1), .rand(r_t39), .z_share0(d4_t39_s0), .z_share1(d4_t39_s1));
  assign r_t39 = stage4_share0[6];
  and_module u_and_t40_d4 (.clk(clk), .x_share0(d3_P0_20_s0), .x_share1(d3_P0_20_s1), .y_share0(d3_G2_19_s0), .y_share1(d3_G2_19_s1), .rand(r_t40), .z_share0(d4_t40_s0), .z_share1(d4_t40_s1));
  assign r_t40 = stage4_share0[10];
  and_module u_and_t41_d4 (.clk(clk), .x_share0(d3_P1_21_s0), .x_share1(d3_P1_21_s1), .y_share0(d3_G2_19_s0), .y_share1(d3_G2_19_s1), .rand(r_t41), .z_share0(d4_t41_s0), .z_share1(d4_t41_s1));
  assign r_t41 = stage4_share0[10];
  and_module u_and_t42_d4 (.clk(clk), .x_share0(d3_P2_22_s0), .x_share1(d3_P2_22_s1), .y_share0(d3_G2_19_s0), .y_share1(d3_G2_19_s1), .rand(r_t42), .z_share0(d4_t42_s0), .z_share1(d4_t42_s1));
  assign r_t42 = stage4_share0[11];
  and_module u_and_t43_d4 (.clk(clk), .x_share0(d3_P2_23_s0), .x_share1(d3_P2_23_s1), .y_share0(d3_G2_19_s0), .y_share1(d3_G2_19_s1), .rand(r_t43), .z_share0(d4_t43_s0), .z_share1(d4_t43_s1));
  assign r_t43 = stage4_share0[11];
  and_module u_and_t44_d4 (.clk(clk), .x_share0(d3_P0_28_s0), .x_share1(d3_P0_28_s1), .y_share0(d3_G2_27_s0), .y_share1(d3_G2_27_s1), .rand(r_t44), .z_share0(d4_t44_s0), .z_share1(d4_t44_s1));
  assign r_t44 = stage4_share0[22];
  and_module u_and_t45_d4 (.clk(clk), .x_share0(d3_P1_29_s0), .x_share1(d3_P1_29_s1), .y_share0(d3_G2_27_s0), .y_share1(d3_G2_27_s1), .rand(r_t45), .z_share0(d4_t45_s0), .z_share1(d4_t45_s1));
  assign r_t45 = stage4_share0[24];
  and_module u_and_t46_d4 (.clk(clk), .x_share0(d3_P2_30_s0), .x_share1(d3_P2_30_s1), .y_share0(d3_G2_27_s0), .y_share1(d3_G2_27_s1), .rand(r_t46), .z_share0(d4_t46_s0), .z_share1(d4_t46_s1));
  assign r_t46 = stage4_share0[22];
  and_module u_and_t47_d4 (.clk(clk), .x_share0(d3_P2_31_s0), .x_share1(d3_P2_31_s1), .y_share0(d3_G2_27_s0), .y_share1(d3_G2_27_s1), .rand(r_t47), .z_share0(d4_t47_s0), .z_share1(d4_t47_s1));
  assign r_t47 = stage4_share0[22];
  reg_module u_reg_G0_16_d5 (.clk(clk), .input_share0(d4_G0_16_s0), .input_share1(d4_G0_16_s1), .output_share0(d5_G0_16_s0), .output_share1(d5_G0_16_s1));
  reg_module u_reg_G0_24_d5 (.clk(clk), .input_share0(d4_G0_24_s0), .input_share1(d4_G0_24_s1), .output_share0(d5_G0_24_s0), .output_share1(d5_G0_24_s1));
  reg_module u_reg_G0_8_d5 (.clk(clk), .input_share0(d4_G0_8_s0), .input_share1(d4_G0_8_s1), .output_share0(d5_G0_8_s0), .output_share1(d5_G0_8_s1));
  reg_module u_reg_G1_17_d5 (.clk(clk), .input_share0(d4_G1_17_s0), .input_share1(d4_G1_17_s1), .output_share0(d5_G1_17_s0), .output_share1(d5_G1_17_s1));
  reg_module u_reg_G1_25_d5 (.clk(clk), .input_share0(d4_G1_25_s0), .input_share1(d4_G1_25_s1), .output_share0(d5_G1_25_s0), .output_share1(d5_G1_25_s1));
  reg_module u_reg_G1_9_d5 (.clk(clk), .input_share0(d4_G1_9_s0), .input_share1(d4_G1_9_s1), .output_share0(d5_G1_9_s0), .output_share1(d5_G1_9_s1));
  reg_module u_reg_G2_10_d5 (.clk(clk), .input_share0(d4_G2_10_s0), .input_share1(d4_G2_10_s1), .output_share0(d5_G2_10_s0), .output_share1(d5_G2_10_s1));
  reg_module u_reg_G2_11_d5 (.clk(clk), .input_share0(d4_G2_11_s0), .input_share1(d4_G2_11_s1), .output_share0(d5_G2_11_s0), .output_share1(d5_G2_11_s1));
  reg_module u_reg_G2_18_d5 (.clk(clk), .input_share0(d4_G2_18_s0), .input_share1(d4_G2_18_s1), .output_share0(d5_G2_18_s0), .output_share1(d5_G2_18_s1));
  reg_module u_reg_G2_19_d5 (.clk(clk), .input_share0(d4_G2_19_s0), .input_share1(d4_G2_19_s1), .output_share0(d5_G2_19_s0), .output_share1(d5_G2_19_s1));
  reg_module u_reg_G2_26_d5 (.clk(clk), .input_share0(d4_G2_26_s0), .input_share1(d4_G2_26_s1), .output_share0(d5_G2_26_s0), .output_share1(d5_G2_26_s1));
  reg_module u_reg_G2_27_d5 (.clk(clk), .input_share0(d4_G2_27_s0), .input_share1(d4_G2_27_s1), .output_share0(d5_G2_27_s0), .output_share1(d5_G2_27_s1));
  reg_module u_reg_G3_12_d5 (.clk(clk), .input_share0(d4_G3_12_s0), .input_share1(d4_G3_12_s1), .output_share0(d5_G3_12_s0), .output_share1(d5_G3_12_s1));
  reg_module u_reg_G3_13_d5 (.clk(clk), .input_share0(d4_G3_13_s0), .input_share1(d4_G3_13_s1), .output_share0(d5_G3_13_s0), .output_share1(d5_G3_13_s1));
  reg_module u_reg_G3_14_d5 (.clk(clk), .input_share0(d4_G3_14_s0), .input_share1(d4_G3_14_s1), .output_share0(d5_G3_14_s0), .output_share1(d5_G3_14_s1));
  reg_module u_reg_G3_15_d5 (.clk(clk), .input_share0(d4_G3_15_s0), .input_share1(d4_G3_15_s1), .output_share0(d5_G3_15_s0), .output_share1(d5_G3_15_s1));
  reg_module u_reg_G3_20_d5 (.clk(clk), .input_share0(d4_G3_20_s0), .input_share1(d4_G3_20_s1), .output_share0(d5_G3_20_s0), .output_share1(d5_G3_20_s1));
  reg_module u_reg_G3_21_d5 (.clk(clk), .input_share0(d4_G3_21_s0), .input_share1(d4_G3_21_s1), .output_share0(d5_G3_21_s0), .output_share1(d5_G3_21_s1));
  reg_module u_reg_G3_22_d5 (.clk(clk), .input_share0(d4_G3_22_s0), .input_share1(d4_G3_22_s1), .output_share0(d5_G3_22_s0), .output_share1(d5_G3_22_s1));
  reg_module u_reg_G3_23_d5 (.clk(clk), .input_share0(d4_G3_23_s0), .input_share1(d4_G3_23_s1), .output_share0(d5_G3_23_s0), .output_share1(d5_G3_23_s1));
  reg_module u_reg_G3_28_d5 (.clk(clk), .input_share0(d4_G3_28_s0), .input_share1(d4_G3_28_s1), .output_share0(d5_G3_28_s0), .output_share1(d5_G3_28_s1));
  reg_module u_reg_G3_29_d5 (.clk(clk), .input_share0(d4_G3_29_s0), .input_share1(d4_G3_29_s1), .output_share0(d5_G3_29_s0), .output_share1(d5_G3_29_s1));
  reg_module u_reg_G3_30_d5 (.clk(clk), .input_share0(d4_G3_30_s0), .input_share1(d4_G3_30_s1), .output_share0(d5_G3_30_s0), .output_share1(d5_G3_30_s1));
  reg_module u_reg_G3_31_d5 (.clk(clk), .input_share0(d4_G3_31_s0), .input_share1(d4_G3_31_s1), .output_share0(d5_G3_31_s0), .output_share1(d5_G3_31_s1));
  reg_module u_reg_P0_10_d5 (.clk(clk), .input_share0(d4_P0_10_s0), .input_share1(d4_P0_10_s1), .output_share0(d5_P0_10_s0), .output_share1(d5_P0_10_s1));
  reg_module u_reg_P0_11_d5 (.clk(clk), .input_share0(d4_P0_11_s0), .input_share1(d4_P0_11_s1), .output_share0(d5_P0_11_s0), .output_share1(d5_P0_11_s1));
  reg_module u_reg_P0_12_d5 (.clk(clk), .input_share0(d4_P0_12_s0), .input_share1(d4_P0_12_s1), .output_share0(d5_P0_12_s0), .output_share1(d5_P0_12_s1));
  reg_module u_reg_P0_13_d5 (.clk(clk), .input_share0(d4_P0_13_s0), .input_share1(d4_P0_13_s1), .output_share0(d5_P0_13_s0), .output_share1(d5_P0_13_s1));
  reg_module u_reg_P0_14_d5 (.clk(clk), .input_share0(d4_P0_14_s0), .input_share1(d4_P0_14_s1), .output_share0(d5_P0_14_s0), .output_share1(d5_P0_14_s1));
  reg_module u_reg_P0_15_d5 (.clk(clk), .input_share0(d4_P0_15_s0), .input_share1(d4_P0_15_s1), .output_share0(d5_P0_15_s0), .output_share1(d5_P0_15_s1));
  reg_module u_reg_P0_16_d5 (.clk(clk), .input_share0(d4_P0_16_s0), .input_share1(d4_P0_16_s1), .output_share0(d5_P0_16_s0), .output_share1(d5_P0_16_s1));
  reg_module u_reg_P0_17_d5 (.clk(clk), .input_share0(d4_P0_17_s0), .input_share1(d4_P0_17_s1), .output_share0(d5_P0_17_s0), .output_share1(d5_P0_17_s1));
  reg_module u_reg_P0_18_d5 (.clk(clk), .input_share0(d4_P0_18_s0), .input_share1(d4_P0_18_s1), .output_share0(d5_P0_18_s0), .output_share1(d5_P0_18_s1));
  reg_module u_reg_P0_19_d5 (.clk(clk), .input_share0(d4_P0_19_s0), .input_share1(d4_P0_19_s1), .output_share0(d5_P0_19_s0), .output_share1(d5_P0_19_s1));
  reg_module u_reg_P0_20_d5 (.clk(clk), .input_share0(d4_P0_20_s0), .input_share1(d4_P0_20_s1), .output_share0(d5_P0_20_s0), .output_share1(d5_P0_20_s1));
  reg_module u_reg_P0_21_d5 (.clk(clk), .input_share0(d4_P0_21_s0), .input_share1(d4_P0_21_s1), .output_share0(d5_P0_21_s0), .output_share1(d5_P0_21_s1));
  reg_module u_reg_P0_22_d5 (.clk(clk), .input_share0(d4_P0_22_s0), .input_share1(d4_P0_22_s1), .output_share0(d5_P0_22_s0), .output_share1(d5_P0_22_s1));
  reg_module u_reg_P0_23_d5 (.clk(clk), .input_share0(d4_P0_23_s0), .input_share1(d4_P0_23_s1), .output_share0(d5_P0_23_s0), .output_share1(d5_P0_23_s1));
  reg_module u_reg_P0_24_d5 (.clk(clk), .input_share0(d4_P0_24_s0), .input_share1(d4_P0_24_s1), .output_share0(d5_P0_24_s0), .output_share1(d5_P0_24_s1));
  reg_module u_reg_P0_25_d5 (.clk(clk), .input_share0(d4_P0_25_s0), .input_share1(d4_P0_25_s1), .output_share0(d5_P0_25_s0), .output_share1(d5_P0_25_s1));
  reg_module u_reg_P0_26_d5 (.clk(clk), .input_share0(d4_P0_26_s0), .input_share1(d4_P0_26_s1), .output_share0(d5_P0_26_s0), .output_share1(d5_P0_26_s1));
  reg_module u_reg_P0_27_d5 (.clk(clk), .input_share0(d4_P0_27_s0), .input_share1(d4_P0_27_s1), .output_share0(d5_P0_27_s0), .output_share1(d5_P0_27_s1));
  reg_module u_reg_P0_28_d5 (.clk(clk), .input_share0(d4_P0_28_s0), .input_share1(d4_P0_28_s1), .output_share0(d5_P0_28_s0), .output_share1(d5_P0_28_s1));
  reg_module u_reg_P0_29_d5 (.clk(clk), .input_share0(d4_P0_29_s0), .input_share1(d4_P0_29_s1), .output_share0(d5_P0_29_s0), .output_share1(d5_P0_29_s1));
  reg_module u_reg_P0_30_d5 (.clk(clk), .input_share0(d4_P0_30_s0), .input_share1(d4_P0_30_s1), .output_share0(d5_P0_30_s0), .output_share1(d5_P0_30_s1));
  reg_module u_reg_P0_31_d5 (.clk(clk), .input_share0(d4_P0_31_s0), .input_share1(d4_P0_31_s1), .output_share0(d5_P0_31_s0), .output_share1(d5_P0_31_s1));
  reg_module u_reg_P0_9_d5 (.clk(clk), .input_share0(d4_P0_9_s0), .input_share1(d4_P0_9_s1), .output_share0(d5_P0_9_s0), .output_share1(d5_P0_9_s1));
  reg_module u_reg_P1_17_d5 (.clk(clk), .input_share0(d4_P1_17_s0), .input_share1(d4_P1_17_s1), .output_share0(d5_P1_17_s0), .output_share1(d5_P1_17_s1));
  reg_module u_reg_P2_18_d5 (.clk(clk), .input_share0(d4_P2_18_s0), .input_share1(d4_P2_18_s1), .output_share0(d5_P2_18_s0), .output_share1(d5_P2_18_s1));
  reg_module u_reg_P2_19_d5 (.clk(clk), .input_share0(d4_P2_19_s0), .input_share1(d4_P2_19_s1), .output_share0(d5_P2_19_s0), .output_share1(d5_P2_19_s1));
  reg_module u_reg_P3_20_d5 (.clk(clk), .input_share0(d4_P3_20_s0), .input_share1(d4_P3_20_s1), .output_share0(d5_P3_20_s0), .output_share1(d5_P3_20_s1));
  reg_module u_reg_P3_21_d5 (.clk(clk), .input_share0(d4_P3_21_s0), .input_share1(d4_P3_21_s1), .output_share0(d5_P3_21_s0), .output_share1(d5_P3_21_s1));
  reg_module u_reg_P3_22_d5 (.clk(clk), .input_share0(d4_P3_22_s0), .input_share1(d4_P3_22_s1), .output_share0(d5_P3_22_s0), .output_share1(d5_P3_22_s1));
  reg_module u_reg_P3_23_d5 (.clk(clk), .input_share0(d4_P3_23_s0), .input_share1(d4_P3_23_s1), .output_share0(d5_P3_23_s0), .output_share1(d5_P3_23_s1));
  reg_module u_reg_P4_24_d5 (.clk(clk), .input_share0(d4_P4_24_s0), .input_share1(d4_P4_24_s1), .output_share0(d5_P4_24_s0), .output_share1(d5_P4_24_s1));
  reg_module u_reg_P4_25_d5 (.clk(clk), .input_share0(d4_P4_25_s0), .input_share1(d4_P4_25_s1), .output_share0(d5_P4_25_s0), .output_share1(d5_P4_25_s1));
  reg_module u_reg_P4_26_d5 (.clk(clk), .input_share0(d4_P4_26_s0), .input_share1(d4_P4_26_s1), .output_share0(d5_P4_26_s0), .output_share1(d5_P4_26_s1));
  reg_module u_reg_P4_27_d5 (.clk(clk), .input_share0(d4_P4_27_s0), .input_share1(d4_P4_27_s1), .output_share0(d5_P4_27_s0), .output_share1(d5_P4_27_s1));
  reg_module u_reg_P4_28_d5 (.clk(clk), .input_share0(d4_P4_28_s0), .input_share1(d4_P4_28_s1), .output_share0(d5_P4_28_s0), .output_share1(d5_P4_28_s1));
  reg_module u_reg_P4_29_d5 (.clk(clk), .input_share0(d4_P4_29_s0), .input_share1(d4_P4_29_s1), .output_share0(d5_P4_29_s0), .output_share1(d5_P4_29_s1));
  reg_module u_reg_P4_30_d5 (.clk(clk), .input_share0(d4_P4_30_s0), .input_share1(d4_P4_30_s1), .output_share0(d5_P4_30_s0), .output_share1(d5_P4_30_s1));
  reg_module u_reg_P4_31_d5 (.clk(clk), .input_share0(d4_P4_31_s0), .input_share1(d4_P4_31_s1), .output_share0(d5_P4_31_s0), .output_share1(d5_P4_31_s1));
  xor_module u_xor_G4_10_d5 (.x_share0(d5_t50_s0), .x_share1(d5_t50_s1), .y_share0(d5_G2_10_s0), .y_share1(d5_G2_10_s1), .z_share0(d5_G4_10_s0), .z_share1(d5_G4_10_s1));
  xor_module u_xor_G4_11_d5 (.x_share0(d5_t51_s0), .x_share1(d5_t51_s1), .y_share0(d5_G2_11_s0), .y_share1(d5_G2_11_s1), .z_share0(d5_G4_11_s0), .z_share1(d5_G4_11_s1));
  xor_module u_xor_G4_12_d5 (.x_share0(d5_t52_s0), .x_share1(d5_t52_s1), .y_share0(d5_G3_12_s0), .y_share1(d5_G3_12_s1), .z_share0(d5_G4_12_s0), .z_share1(d5_G4_12_s1));
  xor_module u_xor_G4_13_d5 (.x_share0(d5_t53_s0), .x_share1(d5_t53_s1), .y_share0(d5_G3_13_s0), .y_share1(d5_G3_13_s1), .z_share0(d5_G4_13_s0), .z_share1(d5_G4_13_s1));
  xor_module u_xor_G4_14_d5 (.x_share0(d5_t54_s0), .x_share1(d5_t54_s1), .y_share0(d5_G3_14_s0), .y_share1(d5_G3_14_s1), .z_share0(d5_G4_14_s0), .z_share1(d5_G4_14_s1));
  xor_module u_xor_G4_15_d5 (.x_share0(d5_t55_s0), .x_share1(d5_t55_s1), .y_share0(d5_G3_15_s0), .y_share1(d5_G3_15_s1), .z_share0(d5_G4_15_s0), .z_share1(d5_G4_15_s1));
  xor_module u_xor_G4_24_d5 (.x_share0(d5_t56_s0), .x_share1(d5_t56_s1), .y_share0(d5_G0_24_s0), .y_share1(d5_G0_24_s1), .z_share0(d5_G4_24_s0), .z_share1(d5_G4_24_s1));
  xor_module u_xor_G4_25_d5 (.x_share0(d5_t57_s0), .x_share1(d5_t57_s1), .y_share0(d5_G1_25_s0), .y_share1(d5_G1_25_s1), .z_share0(d5_G4_25_s0), .z_share1(d5_G4_25_s1));
  xor_module u_xor_G4_26_d5 (.x_share0(d5_t58_s0), .x_share1(d5_t58_s1), .y_share0(d5_G2_26_s0), .y_share1(d5_G2_26_s1), .z_share0(d5_G4_26_s0), .z_share1(d5_G4_26_s1));
  xor_module u_xor_G4_27_d5 (.x_share0(d5_t59_s0), .x_share1(d5_t59_s1), .y_share0(d5_G2_27_s0), .y_share1(d5_G2_27_s1), .z_share0(d5_G4_27_s0), .z_share1(d5_G4_27_s1));
  xor_module u_xor_G4_28_d5 (.x_share0(d5_t60_s0), .x_share1(d5_t60_s1), .y_share0(d5_G3_28_s0), .y_share1(d5_G3_28_s1), .z_share0(d5_G4_28_s0), .z_share1(d5_G4_28_s1));
  xor_module u_xor_G4_29_d5 (.x_share0(d5_t61_s0), .x_share1(d5_t61_s1), .y_share0(d5_G3_29_s0), .y_share1(d5_G3_29_s1), .z_share0(d5_G4_29_s0), .z_share1(d5_G4_29_s1));
  xor_module u_xor_G4_30_d5 (.x_share0(d5_t62_s0), .x_share1(d5_t62_s1), .y_share0(d5_G3_30_s0), .y_share1(d5_G3_30_s1), .z_share0(d5_G4_30_s0), .z_share1(d5_G4_30_s1));
  xor_module u_xor_G4_31_d5 (.x_share0(d5_t63_s0), .x_share1(d5_t63_s1), .y_share0(d5_G3_31_s0), .y_share1(d5_G3_31_s1), .z_share0(d5_G4_31_s0), .z_share1(d5_G4_31_s1));
  xor_module u_xor_G4_8_d5 (.x_share0(d5_t48_s0), .x_share1(d5_t48_s1), .y_share0(d5_G0_8_s0), .y_share1(d5_G0_8_s1), .z_share0(d5_G4_8_s0), .z_share1(d5_G4_8_s1));
  xor_module u_xor_G4_9_d5 (.x_share0(d5_t49_s0), .x_share1(d5_t49_s1), .y_share0(d5_G1_9_s0), .y_share1(d5_G1_9_s1), .z_share0(d5_G4_9_s0), .z_share1(d5_G4_9_s1));
  xor_module u_xor_o10_d5 (.x_share0(d5_P0_10_s0), .x_share1(d5_P0_10_s1), .y_share0(d5_G4_9_s0), .y_share1(d5_G4_9_s1), .z_share0(d5_o10_s0), .z_share1(d5_o10_s1));
  xor_module u_xor_o11_d5 (.x_share0(d5_P0_11_s0), .x_share1(d5_P0_11_s1), .y_share0(d5_G4_10_s0), .y_share1(d5_G4_10_s1), .z_share0(d5_o11_s0), .z_share1(d5_o11_s1));
  xor_module u_xor_o12_d5 (.x_share0(d5_P0_12_s0), .x_share1(d5_P0_12_s1), .y_share0(d5_G4_11_s0), .y_share1(d5_G4_11_s1), .z_share0(d5_o12_s0), .z_share1(d5_o12_s1));
  xor_module u_xor_o13_d5 (.x_share0(d5_P0_13_s0), .x_share1(d5_P0_13_s1), .y_share0(d5_G4_12_s0), .y_share1(d5_G4_12_s1), .z_share0(d5_o13_s0), .z_share1(d5_o13_s1));
  xor_module u_xor_o14_d5 (.x_share0(d5_P0_14_s0), .x_share1(d5_P0_14_s1), .y_share0(d5_G4_13_s0), .y_share1(d5_G4_13_s1), .z_share0(d5_o14_s0), .z_share1(d5_o14_s1));
  xor_module u_xor_o15_d5 (.x_share0(d5_P0_15_s0), .x_share1(d5_P0_15_s1), .y_share0(d5_G4_14_s0), .y_share1(d5_G4_14_s1), .z_share0(d5_o15_s0), .z_share1(d5_o15_s1));
  xor_module u_xor_o16_d5 (.x_share0(d5_P0_16_s0), .x_share1(d5_P0_16_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .z_share0(d5_o16_s0), .z_share1(d5_o16_s1));
  xor_module u_xor_o9_d5 (.x_share0(d5_P0_9_s0), .x_share1(d5_P0_9_s1), .y_share0(d5_G4_8_s0), .y_share1(d5_G4_8_s1), .z_share0(d5_o9_s0), .z_share1(d5_o9_s1));
  and_module u_and_t48_d5 (.clk(clk), .x_share0(d4_P0_8_s0), .x_share1(d4_P0_8_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t48), .z_share0(d5_t48_s0), .z_share1(d5_t48_s1));
  assign r_t48 = stage5_share0[1];
  and_module u_and_t49_d5 (.clk(clk), .x_share0(d4_P1_9_s0), .x_share1(d4_P1_9_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t49), .z_share0(d5_t49_s0), .z_share1(d5_t49_s1));
  assign r_t49 = stage5_share0[0];
  and_module u_and_t50_d5 (.clk(clk), .x_share0(d4_P2_10_s0), .x_share1(d4_P2_10_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t50), .z_share0(d5_t50_s0), .z_share1(d5_t50_s1));
  assign r_t50 = stage5_share0[2];
  and_module u_and_t51_d5 (.clk(clk), .x_share0(d4_P2_11_s0), .x_share1(d4_P2_11_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t51), .z_share0(d5_t51_s0), .z_share1(d5_t51_s1));
  assign r_t51 = stage5_share0[0];
  and_module u_and_t52_d5 (.clk(clk), .x_share0(d4_P3_12_s0), .x_share1(d4_P3_12_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t52), .z_share0(d5_t52_s0), .z_share1(d5_t52_s1));
  assign r_t52 = stage5_share0[2];
  and_module u_and_t53_d5 (.clk(clk), .x_share0(d4_P3_13_s0), .x_share1(d4_P3_13_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t53), .z_share0(d5_t53_s0), .z_share1(d5_t53_s1));
  assign r_t53 = stage5_share0[4];
  and_module u_and_t54_d5 (.clk(clk), .x_share0(d4_P3_14_s0), .x_share1(d4_P3_14_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t54), .z_share0(d5_t54_s0), .z_share1(d5_t54_s1));
  assign r_t54 = stage5_share0[6];
  and_module u_and_t55_d5 (.clk(clk), .x_share0(d4_P3_15_s0), .x_share1(d4_P3_15_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t55), .z_share0(d5_t55_s0), .z_share1(d5_t55_s1));
  assign r_t55 = stage5_share0[7];
  and_module u_and_t56_d5 (.clk(clk), .x_share0(d4_P0_24_s0), .x_share1(d4_P0_24_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t56), .z_share0(d5_t56_s0), .z_share1(d5_t56_s1));
  assign r_t56 = stage5_share0[18];
  and_module u_and_t57_d5 (.clk(clk), .x_share0(d4_P1_25_s0), .x_share1(d4_P1_25_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t57), .z_share0(d5_t57_s0), .z_share1(d5_t57_s1));
  assign r_t57 = stage5_share0[19];
  and_module u_and_t58_d5 (.clk(clk), .x_share0(d4_P2_26_s0), .x_share1(d4_P2_26_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t58), .z_share0(d5_t58_s0), .z_share1(d5_t58_s1));
  assign r_t58 = stage5_share0[18];
  and_module u_and_t59_d5 (.clk(clk), .x_share0(d4_P2_27_s0), .x_share1(d4_P2_27_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t59), .z_share0(d5_t59_s0), .z_share1(d5_t59_s1));
  assign r_t59 = stage5_share0[18];
  and_module u_and_t60_d5 (.clk(clk), .x_share0(d4_P3_28_s0), .x_share1(d4_P3_28_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t60), .z_share0(d5_t60_s0), .z_share1(d5_t60_s1));
  assign r_t60 = stage5_share0[17];
  and_module u_and_t61_d5 (.clk(clk), .x_share0(d4_P3_29_s0), .x_share1(d4_P3_29_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t61), .z_share0(d5_t61_s0), .z_share1(d5_t61_s1));
  assign r_t61 = stage5_share0[17];
  and_module u_and_t62_d5 (.clk(clk), .x_share0(d4_P3_30_s0), .x_share1(d4_P3_30_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t62), .z_share0(d5_t62_s0), .z_share1(d5_t62_s1));
  assign r_t62 = stage5_share0[17];
  and_module u_and_t63_d5 (.clk(clk), .x_share0(d4_P3_31_s0), .x_share1(d4_P3_31_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t63), .z_share0(d5_t63_s0), .z_share1(d5_t63_s1));
  assign r_t63 = stage5_share0[17];
  reg_module u_reg_G0_16_d6 (.clk(clk), .input_share0(d5_G0_16_s0), .input_share1(d5_G0_16_s1), .output_share0(d6_G0_16_s0), .output_share1(d6_G0_16_s1));
  reg_module u_reg_G1_17_d6 (.clk(clk), .input_share0(d5_G1_17_s0), .input_share1(d5_G1_17_s1), .output_share0(d6_G1_17_s0), .output_share1(d6_G1_17_s1));
  reg_module u_reg_G2_18_d6 (.clk(clk), .input_share0(d5_G2_18_s0), .input_share1(d5_G2_18_s1), .output_share0(d6_G2_18_s0), .output_share1(d6_G2_18_s1));
  reg_module u_reg_G2_19_d6 (.clk(clk), .input_share0(d5_G2_19_s0), .input_share1(d5_G2_19_s1), .output_share0(d6_G2_19_s0), .output_share1(d6_G2_19_s1));
  reg_module u_reg_G3_20_d6 (.clk(clk), .input_share0(d5_G3_20_s0), .input_share1(d5_G3_20_s1), .output_share0(d6_G3_20_s0), .output_share1(d6_G3_20_s1));
  reg_module u_reg_G3_21_d6 (.clk(clk), .input_share0(d5_G3_21_s0), .input_share1(d5_G3_21_s1), .output_share0(d6_G3_21_s0), .output_share1(d6_G3_21_s1));
  reg_module u_reg_G3_22_d6 (.clk(clk), .input_share0(d5_G3_22_s0), .input_share1(d5_G3_22_s1), .output_share0(d6_G3_22_s0), .output_share1(d6_G3_22_s1));
  reg_module u_reg_G3_23_d6 (.clk(clk), .input_share0(d5_G3_23_s0), .input_share1(d5_G3_23_s1), .output_share0(d6_G3_23_s0), .output_share1(d6_G3_23_s1));
  reg_module u_reg_G4_24_d6 (.clk(clk), .input_share0(d5_G4_24_s0), .input_share1(d5_G4_24_s1), .output_share0(d6_G4_24_s0), .output_share1(d6_G4_24_s1));
  reg_module u_reg_G4_25_d6 (.clk(clk), .input_share0(d5_G4_25_s0), .input_share1(d5_G4_25_s1), .output_share0(d6_G4_25_s0), .output_share1(d6_G4_25_s1));
  reg_module u_reg_G4_26_d6 (.clk(clk), .input_share0(d5_G4_26_s0), .input_share1(d5_G4_26_s1), .output_share0(d6_G4_26_s0), .output_share1(d6_G4_26_s1));
  reg_module u_reg_G4_27_d6 (.clk(clk), .input_share0(d5_G4_27_s0), .input_share1(d5_G4_27_s1), .output_share0(d6_G4_27_s0), .output_share1(d6_G4_27_s1));
  reg_module u_reg_G4_28_d6 (.clk(clk), .input_share0(d5_G4_28_s0), .input_share1(d5_G4_28_s1), .output_share0(d6_G4_28_s0), .output_share1(d6_G4_28_s1));
  reg_module u_reg_G4_29_d6 (.clk(clk), .input_share0(d5_G4_29_s0), .input_share1(d5_G4_29_s1), .output_share0(d6_G4_29_s0), .output_share1(d6_G4_29_s1));
  reg_module u_reg_G4_30_d6 (.clk(clk), .input_share0(d5_G4_30_s0), .input_share1(d5_G4_30_s1), .output_share0(d6_G4_30_s0), .output_share1(d6_G4_30_s1));
  reg_module u_reg_G4_31_d6 (.clk(clk), .input_share0(d5_G4_31_s0), .input_share1(d5_G4_31_s1), .output_share0(d6_G4_31_s0), .output_share1(d6_G4_31_s1));
  reg_module u_reg_P0_17_d6 (.clk(clk), .input_share0(d5_P0_17_s0), .input_share1(d5_P0_17_s1), .output_share0(d6_P0_17_s0), .output_share1(d6_P0_17_s1));
  reg_module u_reg_P0_18_d6 (.clk(clk), .input_share0(d5_P0_18_s0), .input_share1(d5_P0_18_s1), .output_share0(d6_P0_18_s0), .output_share1(d6_P0_18_s1));
  reg_module u_reg_P0_19_d6 (.clk(clk), .input_share0(d5_P0_19_s0), .input_share1(d5_P0_19_s1), .output_share0(d6_P0_19_s0), .output_share1(d6_P0_19_s1));
  reg_module u_reg_P0_20_d6 (.clk(clk), .input_share0(d5_P0_20_s0), .input_share1(d5_P0_20_s1), .output_share0(d6_P0_20_s0), .output_share1(d6_P0_20_s1));
  reg_module u_reg_P0_21_d6 (.clk(clk), .input_share0(d5_P0_21_s0), .input_share1(d5_P0_21_s1), .output_share0(d6_P0_21_s0), .output_share1(d6_P0_21_s1));
  reg_module u_reg_P0_22_d6 (.clk(clk), .input_share0(d5_P0_22_s0), .input_share1(d5_P0_22_s1), .output_share0(d6_P0_22_s0), .output_share1(d6_P0_22_s1));
  reg_module u_reg_P0_23_d6 (.clk(clk), .input_share0(d5_P0_23_s0), .input_share1(d5_P0_23_s1), .output_share0(d6_P0_23_s0), .output_share1(d6_P0_23_s1));
  reg_module u_reg_P0_24_d6 (.clk(clk), .input_share0(d5_P0_24_s0), .input_share1(d5_P0_24_s1), .output_share0(d6_P0_24_s0), .output_share1(d6_P0_24_s1));
  reg_module u_reg_P0_25_d6 (.clk(clk), .input_share0(d5_P0_25_s0), .input_share1(d5_P0_25_s1), .output_share0(d6_P0_25_s0), .output_share1(d6_P0_25_s1));
  reg_module u_reg_P0_26_d6 (.clk(clk), .input_share0(d5_P0_26_s0), .input_share1(d5_P0_26_s1), .output_share0(d6_P0_26_s0), .output_share1(d6_P0_26_s1));
  reg_module u_reg_P0_27_d6 (.clk(clk), .input_share0(d5_P0_27_s0), .input_share1(d5_P0_27_s1), .output_share0(d6_P0_27_s0), .output_share1(d6_P0_27_s1));
  reg_module u_reg_P0_28_d6 (.clk(clk), .input_share0(d5_P0_28_s0), .input_share1(d5_P0_28_s1), .output_share0(d6_P0_28_s0), .output_share1(d6_P0_28_s1));
  reg_module u_reg_P0_29_d6 (.clk(clk), .input_share0(d5_P0_29_s0), .input_share1(d5_P0_29_s1), .output_share0(d6_P0_29_s0), .output_share1(d6_P0_29_s1));
  reg_module u_reg_P0_30_d6 (.clk(clk), .input_share0(d5_P0_30_s0), .input_share1(d5_P0_30_s1), .output_share0(d6_P0_30_s0), .output_share1(d6_P0_30_s1));
  reg_module u_reg_P0_31_d6 (.clk(clk), .input_share0(d5_P0_31_s0), .input_share1(d5_P0_31_s1), .output_share0(d6_P0_31_s0), .output_share1(d6_P0_31_s1));
  xor_module u_xor_G5_16_d6 (.x_share0(d6_t64_s0), .x_share1(d6_t64_s1), .y_share0(d6_G0_16_s0), .y_share1(d6_G0_16_s1), .z_share0(d6_G5_16_s0), .z_share1(d6_G5_16_s1));
  xor_module u_xor_G5_17_d6 (.x_share0(d6_t65_s0), .x_share1(d6_t65_s1), .y_share0(d6_G1_17_s0), .y_share1(d6_G1_17_s1), .z_share0(d6_G5_17_s0), .z_share1(d6_G5_17_s1));
  xor_module u_xor_G5_18_d6 (.x_share0(d6_t66_s0), .x_share1(d6_t66_s1), .y_share0(d6_G2_18_s0), .y_share1(d6_G2_18_s1), .z_share0(d6_G5_18_s0), .z_share1(d6_G5_18_s1));
  xor_module u_xor_G5_19_d6 (.x_share0(d6_t67_s0), .x_share1(d6_t67_s1), .y_share0(d6_G2_19_s0), .y_share1(d6_G2_19_s1), .z_share0(d6_G5_19_s0), .z_share1(d6_G5_19_s1));
  xor_module u_xor_G5_20_d6 (.x_share0(d6_t68_s0), .x_share1(d6_t68_s1), .y_share0(d6_G3_20_s0), .y_share1(d6_G3_20_s1), .z_share0(d6_G5_20_s0), .z_share1(d6_G5_20_s1));
  xor_module u_xor_G5_21_d6 (.x_share0(d6_t69_s0), .x_share1(d6_t69_s1), .y_share0(d6_G3_21_s0), .y_share1(d6_G3_21_s1), .z_share0(d6_G5_21_s0), .z_share1(d6_G5_21_s1));
  xor_module u_xor_G5_22_d6 (.x_share0(d6_t70_s0), .x_share1(d6_t70_s1), .y_share0(d6_G3_22_s0), .y_share1(d6_G3_22_s1), .z_share0(d6_G5_22_s0), .z_share1(d6_G5_22_s1));
  xor_module u_xor_G5_23_d6 (.x_share0(d6_t71_s0), .x_share1(d6_t71_s1), .y_share0(d6_G3_23_s0), .y_share1(d6_G3_23_s1), .z_share0(d6_G5_23_s0), .z_share1(d6_G5_23_s1));
  xor_module u_xor_G5_24_d6 (.x_share0(d6_t72_s0), .x_share1(d6_t72_s1), .y_share0(d6_G4_24_s0), .y_share1(d6_G4_24_s1), .z_share0(d6_G5_24_s0), .z_share1(d6_G5_24_s1));
  xor_module u_xor_G5_25_d6 (.x_share0(d6_t73_s0), .x_share1(d6_t73_s1), .y_share0(d6_G4_25_s0), .y_share1(d6_G4_25_s1), .z_share0(d6_G5_25_s0), .z_share1(d6_G5_25_s1));
  xor_module u_xor_G5_26_d6 (.x_share0(d6_t74_s0), .x_share1(d6_t74_s1), .y_share0(d6_G4_26_s0), .y_share1(d6_G4_26_s1), .z_share0(d6_G5_26_s0), .z_share1(d6_G5_26_s1));
  xor_module u_xor_G5_27_d6 (.x_share0(d6_t75_s0), .x_share1(d6_t75_s1), .y_share0(d6_G4_27_s0), .y_share1(d6_G4_27_s1), .z_share0(d6_G5_27_s0), .z_share1(d6_G5_27_s1));
  xor_module u_xor_G5_28_d6 (.x_share0(d6_t76_s0), .x_share1(d6_t76_s1), .y_share0(d6_G4_28_s0), .y_share1(d6_G4_28_s1), .z_share0(d6_G5_28_s0), .z_share1(d6_G5_28_s1));
  xor_module u_xor_G5_29_d6 (.x_share0(d6_t77_s0), .x_share1(d6_t77_s1), .y_share0(d6_G4_29_s0), .y_share1(d6_G4_29_s1), .z_share0(d6_G5_29_s0), .z_share1(d6_G5_29_s1));
  xor_module u_xor_G5_30_d6 (.x_share0(d6_t78_s0), .x_share1(d6_t78_s1), .y_share0(d6_G4_30_s0), .y_share1(d6_G4_30_s1), .z_share0(d6_G5_30_s0), .z_share1(d6_G5_30_s1));
  xor_module u_xor_G5_31_d6 (.x_share0(d6_t79_s0), .x_share1(d6_t79_s1), .y_share0(d6_G4_31_s0), .y_share1(d6_G4_31_s1), .z_share0(d6_G5_31_s0), .z_share1(d6_G5_31_s1));
  xor_module u_xor_o17_d6 (.x_share0(d6_P0_17_s0), .x_share1(d6_P0_17_s1), .y_share0(d6_G5_16_s0), .y_share1(d6_G5_16_s1), .z_share0(d6_o17_s0), .z_share1(d6_o17_s1));
  xor_module u_xor_o18_d6 (.x_share0(d6_P0_18_s0), .x_share1(d6_P0_18_s1), .y_share0(d6_G5_17_s0), .y_share1(d6_G5_17_s1), .z_share0(d6_o18_s0), .z_share1(d6_o18_s1));
  xor_module u_xor_o19_d6 (.x_share0(d6_P0_19_s0), .x_share1(d6_P0_19_s1), .y_share0(d6_G5_18_s0), .y_share1(d6_G5_18_s1), .z_share0(d6_o19_s0), .z_share1(d6_o19_s1));
  xor_module u_xor_o20_d6 (.x_share0(d6_P0_20_s0), .x_share1(d6_P0_20_s1), .y_share0(d6_G5_19_s0), .y_share1(d6_G5_19_s1), .z_share0(d6_o20_s0), .z_share1(d6_o20_s1));
  xor_module u_xor_o21_d6 (.x_share0(d6_P0_21_s0), .x_share1(d6_P0_21_s1), .y_share0(d6_G5_20_s0), .y_share1(d6_G5_20_s1), .z_share0(d6_o21_s0), .z_share1(d6_o21_s1));
  xor_module u_xor_o22_d6 (.x_share0(d6_P0_22_s0), .x_share1(d6_P0_22_s1), .y_share0(d6_G5_21_s0), .y_share1(d6_G5_21_s1), .z_share0(d6_o22_s0), .z_share1(d6_o22_s1));
  xor_module u_xor_o23_d6 (.x_share0(d6_P0_23_s0), .x_share1(d6_P0_23_s1), .y_share0(d6_G5_22_s0), .y_share1(d6_G5_22_s1), .z_share0(d6_o23_s0), .z_share1(d6_o23_s1));
  xor_module u_xor_o24_d6 (.x_share0(d6_P0_24_s0), .x_share1(d6_P0_24_s1), .y_share0(d6_G5_23_s0), .y_share1(d6_G5_23_s1), .z_share0(d6_o24_s0), .z_share1(d6_o24_s1));
  xor_module u_xor_o25_d6 (.x_share0(d6_P0_25_s0), .x_share1(d6_P0_25_s1), .y_share0(d6_G5_24_s0), .y_share1(d6_G5_24_s1), .z_share0(d6_o25_s0), .z_share1(d6_o25_s1));
  xor_module u_xor_o26_d6 (.x_share0(d6_P0_26_s0), .x_share1(d6_P0_26_s1), .y_share0(d6_G5_25_s0), .y_share1(d6_G5_25_s1), .z_share0(d6_o26_s0), .z_share1(d6_o26_s1));
  xor_module u_xor_o27_d6 (.x_share0(d6_P0_27_s0), .x_share1(d6_P0_27_s1), .y_share0(d6_G5_26_s0), .y_share1(d6_G5_26_s1), .z_share0(d6_o27_s0), .z_share1(d6_o27_s1));
  xor_module u_xor_o28_d6 (.x_share0(d6_P0_28_s0), .x_share1(d6_P0_28_s1), .y_share0(d6_G5_27_s0), .y_share1(d6_G5_27_s1), .z_share0(d6_o28_s0), .z_share1(d6_o28_s1));
  xor_module u_xor_o29_d6 (.x_share0(d6_P0_29_s0), .x_share1(d6_P0_29_s1), .y_share0(d6_G5_28_s0), .y_share1(d6_G5_28_s1), .z_share0(d6_o29_s0), .z_share1(d6_o29_s1));
  xor_module u_xor_o30_d6 (.x_share0(d6_P0_30_s0), .x_share1(d6_P0_30_s1), .y_share0(d6_G5_29_s0), .y_share1(d6_G5_29_s1), .z_share0(d6_o30_s0), .z_share1(d6_o30_s1));
  xor_module u_xor_o31_d6 (.x_share0(d6_P0_31_s0), .x_share1(d6_P0_31_s1), .y_share0(d6_G5_30_s0), .y_share1(d6_G5_30_s1), .z_share0(d6_o31_s0), .z_share1(d6_o31_s1));
  and_module u_and_t64_d6 (.clk(clk), .x_share0(d5_P0_16_s0), .x_share1(d5_P0_16_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t64), .z_share0(d6_t64_s0), .z_share1(d6_t64_s1));
  assign r_t64 = stage6_share0[14];
  and_module u_and_t65_d6 (.clk(clk), .x_share0(d5_P1_17_s0), .x_share1(d5_P1_17_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t65), .z_share0(d6_t65_s0), .z_share1(d6_t65_s1));
  assign r_t65 = stage6_share0[14];
  and_module u_and_t66_d6 (.clk(clk), .x_share0(d5_P2_18_s0), .x_share1(d5_P2_18_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t66), .z_share0(d6_t66_s0), .z_share1(d6_t66_s1));
  assign r_t66 = stage6_share0[15];
  and_module u_and_t67_d6 (.clk(clk), .x_share0(d5_P2_19_s0), .x_share1(d5_P2_19_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t67), .z_share0(d6_t67_s0), .z_share1(d6_t67_s1));
  assign r_t67 = stage6_share0[14];
  and_module u_and_t68_d6 (.clk(clk), .x_share0(d5_P3_20_s0), .x_share1(d5_P3_20_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t68), .z_share0(d6_t68_s0), .z_share1(d6_t68_s1));
  assign r_t68 = stage6_share0[15];
  and_module u_and_t69_d6 (.clk(clk), .x_share0(d5_P3_21_s0), .x_share1(d5_P3_21_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t69), .z_share0(d6_t69_s0), .z_share1(d6_t69_s1));
  assign r_t69 = stage6_share0[16];
  and_module u_and_t70_d6 (.clk(clk), .x_share0(d5_P3_22_s0), .x_share1(d5_P3_22_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t70), .z_share0(d6_t70_s0), .z_share1(d6_t70_s1));
  assign r_t70 = stage6_share0[16];
  and_module u_and_t71_d6 (.clk(clk), .x_share0(d5_P3_23_s0), .x_share1(d5_P3_23_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t71), .z_share0(d6_t71_s0), .z_share1(d6_t71_s1));
  assign r_t71 = stage6_share0[16];
  and_module u_and_t72_d6 (.clk(clk), .x_share0(d5_P4_24_s0), .x_share1(d5_P4_24_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t72), .z_share0(d6_t72_s0), .z_share1(d6_t72_s1));
  assign r_t72 = stage6_share0[14];
  and_module u_and_t73_d6 (.clk(clk), .x_share0(d5_P4_25_s0), .x_share1(d5_P4_25_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t73), .z_share0(d6_t73_s0), .z_share1(d6_t73_s1));
  assign r_t73 = stage6_share0[14];
  and_module u_and_t74_d6 (.clk(clk), .x_share0(d5_P4_26_s0), .x_share1(d5_P4_26_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t74), .z_share0(d6_t74_s0), .z_share1(d6_t74_s1));
  assign r_t74 = stage6_share0[14];
  and_module u_and_t75_d6 (.clk(clk), .x_share0(d5_P4_27_s0), .x_share1(d5_P4_27_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t75), .z_share0(d6_t75_s0), .z_share1(d6_t75_s1));
  assign r_t75 = stage6_share0[14];
  and_module u_and_t76_d6 (.clk(clk), .x_share0(d5_P4_28_s0), .x_share1(d5_P4_28_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t76), .z_share0(d6_t76_s0), .z_share1(d6_t76_s1));
  assign r_t76 = stage6_share0[14];
  and_module u_and_t77_d6 (.clk(clk), .x_share0(d5_P4_29_s0), .x_share1(d5_P4_29_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t77), .z_share0(d6_t77_s0), .z_share1(d6_t77_s1));
  assign r_t77 = stage6_share0[14];
  and_module u_and_t78_d6 (.clk(clk), .x_share0(d5_P4_30_s0), .x_share1(d5_P4_30_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t78), .z_share0(d6_t78_s0), .z_share1(d6_t78_s1));
  assign r_t78 = stage6_share0[14];
  and_module u_and_t79_d6 (.clk(clk), .x_share0(d5_P4_31_s0), .x_share1(d5_P4_31_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t79), .z_share0(d6_t79_s0), .z_share1(d6_t79_s1));
  assign r_t79 = stage6_share0[14];

  // Output assignments
  assign o_share0[0] = d0_o0_s0;
  assign o_share1[0] = d0_o0_s1;
  assign o_share0[1] = d1_o1_s0;
  assign o_share1[1] = d1_o1_s1;
  assign o_share0[2] = d2_o2_s0;
  assign o_share1[2] = d2_o2_s1;
  assign o_share0[3] = d3_o3_s0;
  assign o_share1[3] = d3_o3_s1;
  assign o_share0[4] = d3_o4_s0;
  assign o_share1[4] = d3_o4_s1;
  assign o_share0[5] = d4_o5_s0;
  assign o_share1[5] = d4_o5_s1;
  assign o_share0[6] = d4_o6_s0;
  assign o_share1[6] = d4_o6_s1;
  assign o_share0[7] = d4_o7_s0;
  assign o_share1[7] = d4_o7_s1;
  assign o_share0[8] = d4_o8_s0;
  assign o_share1[8] = d4_o8_s1;
  assign o_share0[9] = d5_o9_s0;
  assign o_share1[9] = d5_o9_s1;
  assign o_share0[10] = d5_o10_s0;
  assign o_share1[10] = d5_o10_s1;
  assign o_share0[11] = d5_o11_s0;
  assign o_share1[11] = d5_o11_s1;
  assign o_share0[12] = d5_o12_s0;
  assign o_share1[12] = d5_o12_s1;
  assign o_share0[13] = d5_o13_s0;
  assign o_share1[13] = d5_o13_s1;
  assign o_share0[14] = d5_o14_s0;
  assign o_share1[14] = d5_o14_s1;
  assign o_share0[15] = d5_o15_s0;
  assign o_share1[15] = d5_o15_s1;
  assign o_share0[16] = d5_o16_s0;
  assign o_share1[16] = d5_o16_s1;
  assign o_share0[17] = d6_o17_s0;
  assign o_share1[17] = d6_o17_s1;
  assign o_share0[18] = d6_o18_s0;
  assign o_share1[18] = d6_o18_s1;
  assign o_share0[19] = d6_o19_s0;
  assign o_share1[19] = d6_o19_s1;
  assign o_share0[20] = d6_o20_s0;
  assign o_share1[20] = d6_o20_s1;
  assign o_share0[21] = d6_o21_s0;
  assign o_share1[21] = d6_o21_s1;
  assign o_share0[22] = d6_o22_s0;
  assign o_share1[22] = d6_o22_s1;
  assign o_share0[23] = d6_o23_s0;
  assign o_share1[23] = d6_o23_s1;
  assign o_share0[24] = d6_o24_s0;
  assign o_share1[24] = d6_o24_s1;
  assign o_share0[25] = d6_o25_s0;
  assign o_share1[25] = d6_o25_s1;
  assign o_share0[26] = d6_o26_s0;
  assign o_share1[26] = d6_o26_s1;
  assign o_share0[27] = d6_o27_s0;
  assign o_share1[27] = d6_o27_s1;
  assign o_share0[28] = d6_o28_s0;
  assign o_share1[28] = d6_o28_s1;
  assign o_share0[29] = d6_o29_s0;
  assign o_share1[29] = d6_o29_s1;
  assign o_share0[30] = d6_o30_s0;
  assign o_share1[30] = d6_o30_s1;
  assign o_share0[31] = d6_o31_s0;
  assign o_share1[31] = d6_o31_s1;

endmodule
