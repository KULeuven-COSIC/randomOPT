`timescale 1ns / 1ps


module RC3mod_32 (
  input           clk,
  input  [63:0] share0_in,
  input  [63:0] share1_in,
  input  [2:0] rand_bit_share0,
  input  [2:0] rand_bit_share1,
  output [31:0] o_share0,
  output [31:0] o_share1
);

  // Randomness pipeline
  // depth-1 ANDs use rand_bit_share0 directly; deeper ones use these
  wire   [2:0] stage2_share0, stage3_share0, stage4_share0, stage5_share0, stage6_share0, stage7_share0, stage8_share0, stage9_share0, stage10_share0, stage11_share0, stage12_share0, stage13_share0, stage14_share0, stage15_share0, stage16_share0, stage17_share0, stage18_share0, stage19_share0, stage20_share0, stage21_share0, stage22_share0, stage23_share0, stage24_share0, stage25_share0, stage26_share0, stage27_share0, stage28_share0, stage29_share0, stage30_share0, stage31_share0;

  reg_3bits rand_stage1 (.clk(clk), .input_share0(rand_bit_share0), .output_share0(stage2_share0));
  reg_3bits rand_stage2 (.clk(clk), .input_share0(stage2_share0), .output_share0(stage3_share0));
  reg_3bits rand_stage3 (.clk(clk), .input_share0(stage3_share0), .output_share0(stage4_share0));
  reg_3bits rand_stage4 (.clk(clk), .input_share0(stage4_share0), .output_share0(stage5_share0));
  reg_3bits rand_stage5 (.clk(clk), .input_share0(stage5_share0), .output_share0(stage6_share0));
  reg_3bits rand_stage6 (.clk(clk), .input_share0(stage6_share0), .output_share0(stage7_share0));
  reg_3bits rand_stage7 (.clk(clk), .input_share0(stage7_share0), .output_share0(stage8_share0));
  reg_3bits rand_stage8 (.clk(clk), .input_share0(stage8_share0), .output_share0(stage9_share0));
  reg_3bits rand_stage9 (.clk(clk), .input_share0(stage9_share0), .output_share0(stage10_share0));
  reg_3bits rand_stage10 (.clk(clk), .input_share0(stage10_share0), .output_share0(stage11_share0));
  reg_3bits rand_stage11 (.clk(clk), .input_share0(stage11_share0), .output_share0(stage12_share0));
  reg_3bits rand_stage12 (.clk(clk), .input_share0(stage12_share0), .output_share0(stage13_share0));
  reg_3bits rand_stage13 (.clk(clk), .input_share0(stage13_share0), .output_share0(stage14_share0));
  reg_3bits rand_stage14 (.clk(clk), .input_share0(stage14_share0), .output_share0(stage15_share0));
  reg_3bits rand_stage15 (.clk(clk), .input_share0(stage15_share0), .output_share0(stage16_share0));
  reg_3bits rand_stage16 (.clk(clk), .input_share0(stage16_share0), .output_share0(stage17_share0));
  reg_3bits rand_stage17 (.clk(clk), .input_share0(stage17_share0), .output_share0(stage18_share0));
  reg_3bits rand_stage18 (.clk(clk), .input_share0(stage18_share0), .output_share0(stage19_share0));
  reg_3bits rand_stage19 (.clk(clk), .input_share0(stage19_share0), .output_share0(stage20_share0));
  reg_3bits rand_stage20 (.clk(clk), .input_share0(stage20_share0), .output_share0(stage21_share0));
  reg_3bits rand_stage21 (.clk(clk), .input_share0(stage21_share0), .output_share0(stage22_share0));
  reg_3bits rand_stage22 (.clk(clk), .input_share0(stage22_share0), .output_share0(stage23_share0));
  reg_3bits rand_stage23 (.clk(clk), .input_share0(stage23_share0), .output_share0(stage24_share0));
  reg_3bits rand_stage24 (.clk(clk), .input_share0(stage24_share0), .output_share0(stage25_share0));
  reg_3bits rand_stage25 (.clk(clk), .input_share0(stage25_share0), .output_share0(stage26_share0));
  reg_3bits rand_stage26 (.clk(clk), .input_share0(stage26_share0), .output_share0(stage27_share0));
  reg_3bits rand_stage27 (.clk(clk), .input_share0(stage27_share0), .output_share0(stage28_share0));
  reg_3bits rand_stage28 (.clk(clk), .input_share0(stage28_share0), .output_share0(stage29_share0));
  reg_3bits rand_stage29 (.clk(clk), .input_share0(stage29_share0), .output_share0(stage30_share0));
  reg_3bits rand_stage30 (.clk(clk), .input_share0(stage30_share0), .output_share0(stage31_share0));

  xor_module u_xor_o0_d0 (.x_share0(share0_in[0]), .x_share1(share1_in[0]), .y_share0(share0_in[32]), .y_share1(share1_in[32]), .z_share0(d0_o0_s0), .z_share1(d0_o0_s1));
  xor_module u_xor_t0_1_d0 (.x_share0(share0_in[1]), .x_share1(share1_in[1]), .y_share0(share0_in[33]), .y_share1(share1_in[33]), .z_share0(d0_t0_1_s0), .z_share1(d0_t0_1_s1));
  xor_module u_xor_t0_10_d0 (.x_share0(share0_in[10]), .x_share1(share1_in[10]), .y_share0(share0_in[42]), .y_share1(share1_in[42]), .z_share0(d0_t0_10_s0), .z_share1(d0_t0_10_s1));
  xor_module u_xor_t0_11_d0 (.x_share0(share0_in[11]), .x_share1(share1_in[11]), .y_share0(share0_in[43]), .y_share1(share1_in[43]), .z_share0(d0_t0_11_s0), .z_share1(d0_t0_11_s1));
  xor_module u_xor_t0_12_d0 (.x_share0(share0_in[12]), .x_share1(share1_in[12]), .y_share0(share0_in[44]), .y_share1(share1_in[44]), .z_share0(d0_t0_12_s0), .z_share1(d0_t0_12_s1));
  xor_module u_xor_t0_13_d0 (.x_share0(share0_in[13]), .x_share1(share1_in[13]), .y_share0(share0_in[45]), .y_share1(share1_in[45]), .z_share0(d0_t0_13_s0), .z_share1(d0_t0_13_s1));
  xor_module u_xor_t0_14_d0 (.x_share0(share0_in[14]), .x_share1(share1_in[14]), .y_share0(share0_in[46]), .y_share1(share1_in[46]), .z_share0(d0_t0_14_s0), .z_share1(d0_t0_14_s1));
  xor_module u_xor_t0_15_d0 (.x_share0(share0_in[15]), .x_share1(share1_in[15]), .y_share0(share0_in[47]), .y_share1(share1_in[47]), .z_share0(d0_t0_15_s0), .z_share1(d0_t0_15_s1));
  xor_module u_xor_t0_16_d0 (.x_share0(share0_in[16]), .x_share1(share1_in[16]), .y_share0(share0_in[48]), .y_share1(share1_in[48]), .z_share0(d0_t0_16_s0), .z_share1(d0_t0_16_s1));
  xor_module u_xor_t0_17_d0 (.x_share0(share0_in[17]), .x_share1(share1_in[17]), .y_share0(share0_in[49]), .y_share1(share1_in[49]), .z_share0(d0_t0_17_s0), .z_share1(d0_t0_17_s1));
  xor_module u_xor_t0_18_d0 (.x_share0(share0_in[18]), .x_share1(share1_in[18]), .y_share0(share0_in[50]), .y_share1(share1_in[50]), .z_share0(d0_t0_18_s0), .z_share1(d0_t0_18_s1));
  xor_module u_xor_t0_19_d0 (.x_share0(share0_in[19]), .x_share1(share1_in[19]), .y_share0(share0_in[51]), .y_share1(share1_in[51]), .z_share0(d0_t0_19_s0), .z_share1(d0_t0_19_s1));
  xor_module u_xor_t0_2_d0 (.x_share0(share0_in[2]), .x_share1(share1_in[2]), .y_share0(share0_in[34]), .y_share1(share1_in[34]), .z_share0(d0_t0_2_s0), .z_share1(d0_t0_2_s1));
  xor_module u_xor_t0_20_d0 (.x_share0(share0_in[20]), .x_share1(share1_in[20]), .y_share0(share0_in[52]), .y_share1(share1_in[52]), .z_share0(d0_t0_20_s0), .z_share1(d0_t0_20_s1));
  xor_module u_xor_t0_21_d0 (.x_share0(share0_in[21]), .x_share1(share1_in[21]), .y_share0(share0_in[53]), .y_share1(share1_in[53]), .z_share0(d0_t0_21_s0), .z_share1(d0_t0_21_s1));
  xor_module u_xor_t0_22_d0 (.x_share0(share0_in[22]), .x_share1(share1_in[22]), .y_share0(share0_in[54]), .y_share1(share1_in[54]), .z_share0(d0_t0_22_s0), .z_share1(d0_t0_22_s1));
  xor_module u_xor_t0_23_d0 (.x_share0(share0_in[23]), .x_share1(share1_in[23]), .y_share0(share0_in[55]), .y_share1(share1_in[55]), .z_share0(d0_t0_23_s0), .z_share1(d0_t0_23_s1));
  xor_module u_xor_t0_24_d0 (.x_share0(share0_in[24]), .x_share1(share1_in[24]), .y_share0(share0_in[56]), .y_share1(share1_in[56]), .z_share0(d0_t0_24_s0), .z_share1(d0_t0_24_s1));
  xor_module u_xor_t0_25_d0 (.x_share0(share0_in[25]), .x_share1(share1_in[25]), .y_share0(share0_in[57]), .y_share1(share1_in[57]), .z_share0(d0_t0_25_s0), .z_share1(d0_t0_25_s1));
  xor_module u_xor_t0_26_d0 (.x_share0(share0_in[26]), .x_share1(share1_in[26]), .y_share0(share0_in[58]), .y_share1(share1_in[58]), .z_share0(d0_t0_26_s0), .z_share1(d0_t0_26_s1));
  xor_module u_xor_t0_27_d0 (.x_share0(share0_in[27]), .x_share1(share1_in[27]), .y_share0(share0_in[59]), .y_share1(share1_in[59]), .z_share0(d0_t0_27_s0), .z_share1(d0_t0_27_s1));
  xor_module u_xor_t0_28_d0 (.x_share0(share0_in[28]), .x_share1(share1_in[28]), .y_share0(share0_in[60]), .y_share1(share1_in[60]), .z_share0(d0_t0_28_s0), .z_share1(d0_t0_28_s1));
  xor_module u_xor_t0_29_d0 (.x_share0(share0_in[29]), .x_share1(share1_in[29]), .y_share0(share0_in[61]), .y_share1(share1_in[61]), .z_share0(d0_t0_29_s0), .z_share1(d0_t0_29_s1));
  xor_module u_xor_t0_3_d0 (.x_share0(share0_in[3]), .x_share1(share1_in[3]), .y_share0(share0_in[35]), .y_share1(share1_in[35]), .z_share0(d0_t0_3_s0), .z_share1(d0_t0_3_s1));
  xor_module u_xor_t0_30_d0 (.x_share0(share0_in[30]), .x_share1(share1_in[30]), .y_share0(share0_in[62]), .y_share1(share1_in[62]), .z_share0(d0_t0_30_s0), .z_share1(d0_t0_30_s1));
  xor_module u_xor_t0_31_d0 (.x_share0(share0_in[31]), .x_share1(share1_in[31]), .y_share0(share0_in[63]), .y_share1(share1_in[63]), .z_share0(d0_t0_31_s0), .z_share1(d0_t0_31_s1));
  xor_module u_xor_t0_4_d0 (.x_share0(share0_in[4]), .x_share1(share1_in[4]), .y_share0(share0_in[36]), .y_share1(share1_in[36]), .z_share0(d0_t0_4_s0), .z_share1(d0_t0_4_s1));
  xor_module u_xor_t0_5_d0 (.x_share0(share0_in[5]), .x_share1(share1_in[5]), .y_share0(share0_in[37]), .y_share1(share1_in[37]), .z_share0(d0_t0_5_s0), .z_share1(d0_t0_5_s1));
  xor_module u_xor_t0_6_d0 (.x_share0(share0_in[6]), .x_share1(share1_in[6]), .y_share0(share0_in[38]), .y_share1(share1_in[38]), .z_share0(d0_t0_6_s0), .z_share1(d0_t0_6_s1));
  xor_module u_xor_t0_7_d0 (.x_share0(share0_in[7]), .x_share1(share1_in[7]), .y_share0(share0_in[39]), .y_share1(share1_in[39]), .z_share0(d0_t0_7_s0), .z_share1(d0_t0_7_s1));
  xor_module u_xor_t0_8_d0 (.x_share0(share0_in[8]), .x_share1(share1_in[8]), .y_share0(share0_in[40]), .y_share1(share1_in[40]), .z_share0(d0_t0_8_s0), .z_share1(d0_t0_8_s1));
  xor_module u_xor_t0_9_d0 (.x_share0(share0_in[9]), .x_share1(share1_in[9]), .y_share0(share0_in[41]), .y_share1(share1_in[41]), .z_share0(d0_t0_9_s0), .z_share1(d0_t0_9_s1));
  reg_module u_reg_i1_d1 (.clk(clk), .input_share0(share0_in[1]), .input_share1(share1_in[1]), .output_share0(d1_i1_s0), .output_share1(d1_i1_s1));
  reg_module u_reg_i10_d1 (.clk(clk), .input_share0(share0_in[10]), .input_share1(share1_in[10]), .output_share0(d1_i10_s0), .output_share1(d1_i10_s1));
  reg_module u_reg_i11_d1 (.clk(clk), .input_share0(share0_in[11]), .input_share1(share1_in[11]), .output_share0(d1_i11_s0), .output_share1(d1_i11_s1));
  reg_module u_reg_i12_d1 (.clk(clk), .input_share0(share0_in[12]), .input_share1(share1_in[12]), .output_share0(d1_i12_s0), .output_share1(d1_i12_s1));
  reg_module u_reg_i13_d1 (.clk(clk), .input_share0(share0_in[13]), .input_share1(share1_in[13]), .output_share0(d1_i13_s0), .output_share1(d1_i13_s1));
  reg_module u_reg_i14_d1 (.clk(clk), .input_share0(share0_in[14]), .input_share1(share1_in[14]), .output_share0(d1_i14_s0), .output_share1(d1_i14_s1));
  reg_module u_reg_i15_d1 (.clk(clk), .input_share0(share0_in[15]), .input_share1(share1_in[15]), .output_share0(d1_i15_s0), .output_share1(d1_i15_s1));
  reg_module u_reg_i16_d1 (.clk(clk), .input_share0(share0_in[16]), .input_share1(share1_in[16]), .output_share0(d1_i16_s0), .output_share1(d1_i16_s1));
  reg_module u_reg_i17_d1 (.clk(clk), .input_share0(share0_in[17]), .input_share1(share1_in[17]), .output_share0(d1_i17_s0), .output_share1(d1_i17_s1));
  reg_module u_reg_i18_d1 (.clk(clk), .input_share0(share0_in[18]), .input_share1(share1_in[18]), .output_share0(d1_i18_s0), .output_share1(d1_i18_s1));
  reg_module u_reg_i19_d1 (.clk(clk), .input_share0(share0_in[19]), .input_share1(share1_in[19]), .output_share0(d1_i19_s0), .output_share1(d1_i19_s1));
  reg_module u_reg_i2_d1 (.clk(clk), .input_share0(share0_in[2]), .input_share1(share1_in[2]), .output_share0(d1_i2_s0), .output_share1(d1_i2_s1));
  reg_module u_reg_i20_d1 (.clk(clk), .input_share0(share0_in[20]), .input_share1(share1_in[20]), .output_share0(d1_i20_s0), .output_share1(d1_i20_s1));
  reg_module u_reg_i21_d1 (.clk(clk), .input_share0(share0_in[21]), .input_share1(share1_in[21]), .output_share0(d1_i21_s0), .output_share1(d1_i21_s1));
  reg_module u_reg_i22_d1 (.clk(clk), .input_share0(share0_in[22]), .input_share1(share1_in[22]), .output_share0(d1_i22_s0), .output_share1(d1_i22_s1));
  reg_module u_reg_i23_d1 (.clk(clk), .input_share0(share0_in[23]), .input_share1(share1_in[23]), .output_share0(d1_i23_s0), .output_share1(d1_i23_s1));
  reg_module u_reg_i24_d1 (.clk(clk), .input_share0(share0_in[24]), .input_share1(share1_in[24]), .output_share0(d1_i24_s0), .output_share1(d1_i24_s1));
  reg_module u_reg_i25_d1 (.clk(clk), .input_share0(share0_in[25]), .input_share1(share1_in[25]), .output_share0(d1_i25_s0), .output_share1(d1_i25_s1));
  reg_module u_reg_i26_d1 (.clk(clk), .input_share0(share0_in[26]), .input_share1(share1_in[26]), .output_share0(d1_i26_s0), .output_share1(d1_i26_s1));
  reg_module u_reg_i27_d1 (.clk(clk), .input_share0(share0_in[27]), .input_share1(share1_in[27]), .output_share0(d1_i27_s0), .output_share1(d1_i27_s1));
  reg_module u_reg_i28_d1 (.clk(clk), .input_share0(share0_in[28]), .input_share1(share1_in[28]), .output_share0(d1_i28_s0), .output_share1(d1_i28_s1));
  reg_module u_reg_i29_d1 (.clk(clk), .input_share0(share0_in[29]), .input_share1(share1_in[29]), .output_share0(d1_i29_s0), .output_share1(d1_i29_s1));
  reg_module u_reg_i3_d1 (.clk(clk), .input_share0(share0_in[3]), .input_share1(share1_in[3]), .output_share0(d1_i3_s0), .output_share1(d1_i3_s1));
  reg_module u_reg_i30_d1 (.clk(clk), .input_share0(share0_in[30]), .input_share1(share1_in[30]), .output_share0(d1_i30_s0), .output_share1(d1_i30_s1));
  reg_module u_reg_i4_d1 (.clk(clk), .input_share0(share0_in[4]), .input_share1(share1_in[4]), .output_share0(d1_i4_s0), .output_share1(d1_i4_s1));
  reg_module u_reg_i5_d1 (.clk(clk), .input_share0(share0_in[5]), .input_share1(share1_in[5]), .output_share0(d1_i5_s0), .output_share1(d1_i5_s1));
  reg_module u_reg_i6_d1 (.clk(clk), .input_share0(share0_in[6]), .input_share1(share1_in[6]), .output_share0(d1_i6_s0), .output_share1(d1_i6_s1));
  reg_module u_reg_i7_d1 (.clk(clk), .input_share0(share0_in[7]), .input_share1(share1_in[7]), .output_share0(d1_i7_s0), .output_share1(d1_i7_s1));
  reg_module u_reg_i8_d1 (.clk(clk), .input_share0(share0_in[8]), .input_share1(share1_in[8]), .output_share0(d1_i8_s0), .output_share1(d1_i8_s1));
  reg_module u_reg_i9_d1 (.clk(clk), .input_share0(share0_in[9]), .input_share1(share1_in[9]), .output_share0(d1_i9_s0), .output_share1(d1_i9_s1));
  reg_module u_reg_t0_1_d1 (.clk(clk), .input_share0(d0_t0_1_s0), .input_share1(d0_t0_1_s1), .output_share0(d1_t0_1_s0), .output_share1(d1_t0_1_s1));
  reg_module u_reg_t0_10_d1 (.clk(clk), .input_share0(d0_t0_10_s0), .input_share1(d0_t0_10_s1), .output_share0(d1_t0_10_s0), .output_share1(d1_t0_10_s1));
  reg_module u_reg_t0_11_d1 (.clk(clk), .input_share0(d0_t0_11_s0), .input_share1(d0_t0_11_s1), .output_share0(d1_t0_11_s0), .output_share1(d1_t0_11_s1));
  reg_module u_reg_t0_12_d1 (.clk(clk), .input_share0(d0_t0_12_s0), .input_share1(d0_t0_12_s1), .output_share0(d1_t0_12_s0), .output_share1(d1_t0_12_s1));
  reg_module u_reg_t0_13_d1 (.clk(clk), .input_share0(d0_t0_13_s0), .input_share1(d0_t0_13_s1), .output_share0(d1_t0_13_s0), .output_share1(d1_t0_13_s1));
  reg_module u_reg_t0_14_d1 (.clk(clk), .input_share0(d0_t0_14_s0), .input_share1(d0_t0_14_s1), .output_share0(d1_t0_14_s0), .output_share1(d1_t0_14_s1));
  reg_module u_reg_t0_15_d1 (.clk(clk), .input_share0(d0_t0_15_s0), .input_share1(d0_t0_15_s1), .output_share0(d1_t0_15_s0), .output_share1(d1_t0_15_s1));
  reg_module u_reg_t0_16_d1 (.clk(clk), .input_share0(d0_t0_16_s0), .input_share1(d0_t0_16_s1), .output_share0(d1_t0_16_s0), .output_share1(d1_t0_16_s1));
  reg_module u_reg_t0_17_d1 (.clk(clk), .input_share0(d0_t0_17_s0), .input_share1(d0_t0_17_s1), .output_share0(d1_t0_17_s0), .output_share1(d1_t0_17_s1));
  reg_module u_reg_t0_18_d1 (.clk(clk), .input_share0(d0_t0_18_s0), .input_share1(d0_t0_18_s1), .output_share0(d1_t0_18_s0), .output_share1(d1_t0_18_s1));
  reg_module u_reg_t0_19_d1 (.clk(clk), .input_share0(d0_t0_19_s0), .input_share1(d0_t0_19_s1), .output_share0(d1_t0_19_s0), .output_share1(d1_t0_19_s1));
  reg_module u_reg_t0_2_d1 (.clk(clk), .input_share0(d0_t0_2_s0), .input_share1(d0_t0_2_s1), .output_share0(d1_t0_2_s0), .output_share1(d1_t0_2_s1));
  reg_module u_reg_t0_20_d1 (.clk(clk), .input_share0(d0_t0_20_s0), .input_share1(d0_t0_20_s1), .output_share0(d1_t0_20_s0), .output_share1(d1_t0_20_s1));
  reg_module u_reg_t0_21_d1 (.clk(clk), .input_share0(d0_t0_21_s0), .input_share1(d0_t0_21_s1), .output_share0(d1_t0_21_s0), .output_share1(d1_t0_21_s1));
  reg_module u_reg_t0_22_d1 (.clk(clk), .input_share0(d0_t0_22_s0), .input_share1(d0_t0_22_s1), .output_share0(d1_t0_22_s0), .output_share1(d1_t0_22_s1));
  reg_module u_reg_t0_23_d1 (.clk(clk), .input_share0(d0_t0_23_s0), .input_share1(d0_t0_23_s1), .output_share0(d1_t0_23_s0), .output_share1(d1_t0_23_s1));
  reg_module u_reg_t0_24_d1 (.clk(clk), .input_share0(d0_t0_24_s0), .input_share1(d0_t0_24_s1), .output_share0(d1_t0_24_s0), .output_share1(d1_t0_24_s1));
  reg_module u_reg_t0_25_d1 (.clk(clk), .input_share0(d0_t0_25_s0), .input_share1(d0_t0_25_s1), .output_share0(d1_t0_25_s0), .output_share1(d1_t0_25_s1));
  reg_module u_reg_t0_26_d1 (.clk(clk), .input_share0(d0_t0_26_s0), .input_share1(d0_t0_26_s1), .output_share0(d1_t0_26_s0), .output_share1(d1_t0_26_s1));
  reg_module u_reg_t0_27_d1 (.clk(clk), .input_share0(d0_t0_27_s0), .input_share1(d0_t0_27_s1), .output_share0(d1_t0_27_s0), .output_share1(d1_t0_27_s1));
  reg_module u_reg_t0_28_d1 (.clk(clk), .input_share0(d0_t0_28_s0), .input_share1(d0_t0_28_s1), .output_share0(d1_t0_28_s0), .output_share1(d1_t0_28_s1));
  reg_module u_reg_t0_29_d1 (.clk(clk), .input_share0(d0_t0_29_s0), .input_share1(d0_t0_29_s1), .output_share0(d1_t0_29_s0), .output_share1(d1_t0_29_s1));
  reg_module u_reg_t0_3_d1 (.clk(clk), .input_share0(d0_t0_3_s0), .input_share1(d0_t0_3_s1), .output_share0(d1_t0_3_s0), .output_share1(d1_t0_3_s1));
  reg_module u_reg_t0_30_d1 (.clk(clk), .input_share0(d0_t0_30_s0), .input_share1(d0_t0_30_s1), .output_share0(d1_t0_30_s0), .output_share1(d1_t0_30_s1));
  reg_module u_reg_t0_31_d1 (.clk(clk), .input_share0(d0_t0_31_s0), .input_share1(d0_t0_31_s1), .output_share0(d1_t0_31_s0), .output_share1(d1_t0_31_s1));
  reg_module u_reg_t0_4_d1 (.clk(clk), .input_share0(d0_t0_4_s0), .input_share1(d0_t0_4_s1), .output_share0(d1_t0_4_s0), .output_share1(d1_t0_4_s1));
  reg_module u_reg_t0_5_d1 (.clk(clk), .input_share0(d0_t0_5_s0), .input_share1(d0_t0_5_s1), .output_share0(d1_t0_5_s0), .output_share1(d1_t0_5_s1));
  reg_module u_reg_t0_6_d1 (.clk(clk), .input_share0(d0_t0_6_s0), .input_share1(d0_t0_6_s1), .output_share0(d1_t0_6_s0), .output_share1(d1_t0_6_s1));
  reg_module u_reg_t0_7_d1 (.clk(clk), .input_share0(d0_t0_7_s0), .input_share1(d0_t0_7_s1), .output_share0(d1_t0_7_s0), .output_share1(d1_t0_7_s1));
  reg_module u_reg_t0_8_d1 (.clk(clk), .input_share0(d0_t0_8_s0), .input_share1(d0_t0_8_s1), .output_share0(d1_t0_8_s0), .output_share1(d1_t0_8_s1));
  reg_module u_reg_t0_9_d1 (.clk(clk), .input_share0(d0_t0_9_s0), .input_share1(d0_t0_9_s1), .output_share0(d1_t0_9_s0), .output_share1(d1_t0_9_s1));
  and_module u_and_c1_d1 (.clk(clk), .x_share0(share0_in[0]), .x_share1(share1_in[0]), .y_share0(share0_in[32]), .y_share1(share1_in[32]), .rand(r_c1), .z_share0(d1_c1_s0), .z_share1(d1_c1_s1));
  assign r_c1 = rand_bit_share0[1];
  xor_module u_xor_o1_d1 (.x_share0(d1_t0_1_s0), .x_share1(d1_t0_1_s1), .y_share0(d1_c1_s0), .y_share1(d1_c1_s1), .z_share0(d1_o1_s0), .z_share1(d1_o1_s1));
  xor_module u_xor_t1_1_d1 (.x_share0(d1_i1_s0), .x_share1(d1_i1_s1), .y_share0(d1_c1_s0), .y_share1(d1_c1_s1), .z_share0(d1_t1_1_s0), .z_share1(d1_t1_1_s1));
  reg_module u_reg_i1_d2 (.clk(clk), .input_share0(d1_i1_s0), .input_share1(d1_i1_s1), .output_share0(d2_i1_s0), .output_share1(d2_i1_s1));
  reg_module u_reg_i10_d2 (.clk(clk), .input_share0(d1_i10_s0), .input_share1(d1_i10_s1), .output_share0(d2_i10_s0), .output_share1(d2_i10_s1));
  reg_module u_reg_i11_d2 (.clk(clk), .input_share0(d1_i11_s0), .input_share1(d1_i11_s1), .output_share0(d2_i11_s0), .output_share1(d2_i11_s1));
  reg_module u_reg_i12_d2 (.clk(clk), .input_share0(d1_i12_s0), .input_share1(d1_i12_s1), .output_share0(d2_i12_s0), .output_share1(d2_i12_s1));
  reg_module u_reg_i13_d2 (.clk(clk), .input_share0(d1_i13_s0), .input_share1(d1_i13_s1), .output_share0(d2_i13_s0), .output_share1(d2_i13_s1));
  reg_module u_reg_i14_d2 (.clk(clk), .input_share0(d1_i14_s0), .input_share1(d1_i14_s1), .output_share0(d2_i14_s0), .output_share1(d2_i14_s1));
  reg_module u_reg_i15_d2 (.clk(clk), .input_share0(d1_i15_s0), .input_share1(d1_i15_s1), .output_share0(d2_i15_s0), .output_share1(d2_i15_s1));
  reg_module u_reg_i16_d2 (.clk(clk), .input_share0(d1_i16_s0), .input_share1(d1_i16_s1), .output_share0(d2_i16_s0), .output_share1(d2_i16_s1));
  reg_module u_reg_i17_d2 (.clk(clk), .input_share0(d1_i17_s0), .input_share1(d1_i17_s1), .output_share0(d2_i17_s0), .output_share1(d2_i17_s1));
  reg_module u_reg_i18_d2 (.clk(clk), .input_share0(d1_i18_s0), .input_share1(d1_i18_s1), .output_share0(d2_i18_s0), .output_share1(d2_i18_s1));
  reg_module u_reg_i19_d2 (.clk(clk), .input_share0(d1_i19_s0), .input_share1(d1_i19_s1), .output_share0(d2_i19_s0), .output_share1(d2_i19_s1));
  reg_module u_reg_i2_d2 (.clk(clk), .input_share0(d1_i2_s0), .input_share1(d1_i2_s1), .output_share0(d2_i2_s0), .output_share1(d2_i2_s1));
  reg_module u_reg_i20_d2 (.clk(clk), .input_share0(d1_i20_s0), .input_share1(d1_i20_s1), .output_share0(d2_i20_s0), .output_share1(d2_i20_s1));
  reg_module u_reg_i21_d2 (.clk(clk), .input_share0(d1_i21_s0), .input_share1(d1_i21_s1), .output_share0(d2_i21_s0), .output_share1(d2_i21_s1));
  reg_module u_reg_i22_d2 (.clk(clk), .input_share0(d1_i22_s0), .input_share1(d1_i22_s1), .output_share0(d2_i22_s0), .output_share1(d2_i22_s1));
  reg_module u_reg_i23_d2 (.clk(clk), .input_share0(d1_i23_s0), .input_share1(d1_i23_s1), .output_share0(d2_i23_s0), .output_share1(d2_i23_s1));
  reg_module u_reg_i24_d2 (.clk(clk), .input_share0(d1_i24_s0), .input_share1(d1_i24_s1), .output_share0(d2_i24_s0), .output_share1(d2_i24_s1));
  reg_module u_reg_i25_d2 (.clk(clk), .input_share0(d1_i25_s0), .input_share1(d1_i25_s1), .output_share0(d2_i25_s0), .output_share1(d2_i25_s1));
  reg_module u_reg_i26_d2 (.clk(clk), .input_share0(d1_i26_s0), .input_share1(d1_i26_s1), .output_share0(d2_i26_s0), .output_share1(d2_i26_s1));
  reg_module u_reg_i27_d2 (.clk(clk), .input_share0(d1_i27_s0), .input_share1(d1_i27_s1), .output_share0(d2_i27_s0), .output_share1(d2_i27_s1));
  reg_module u_reg_i28_d2 (.clk(clk), .input_share0(d1_i28_s0), .input_share1(d1_i28_s1), .output_share0(d2_i28_s0), .output_share1(d2_i28_s1));
  reg_module u_reg_i29_d2 (.clk(clk), .input_share0(d1_i29_s0), .input_share1(d1_i29_s1), .output_share0(d2_i29_s0), .output_share1(d2_i29_s1));
  reg_module u_reg_i3_d2 (.clk(clk), .input_share0(d1_i3_s0), .input_share1(d1_i3_s1), .output_share0(d2_i3_s0), .output_share1(d2_i3_s1));
  reg_module u_reg_i30_d2 (.clk(clk), .input_share0(d1_i30_s0), .input_share1(d1_i30_s1), .output_share0(d2_i30_s0), .output_share1(d2_i30_s1));
  reg_module u_reg_i4_d2 (.clk(clk), .input_share0(d1_i4_s0), .input_share1(d1_i4_s1), .output_share0(d2_i4_s0), .output_share1(d2_i4_s1));
  reg_module u_reg_i5_d2 (.clk(clk), .input_share0(d1_i5_s0), .input_share1(d1_i5_s1), .output_share0(d2_i5_s0), .output_share1(d2_i5_s1));
  reg_module u_reg_i6_d2 (.clk(clk), .input_share0(d1_i6_s0), .input_share1(d1_i6_s1), .output_share0(d2_i6_s0), .output_share1(d2_i6_s1));
  reg_module u_reg_i7_d2 (.clk(clk), .input_share0(d1_i7_s0), .input_share1(d1_i7_s1), .output_share0(d2_i7_s0), .output_share1(d2_i7_s1));
  reg_module u_reg_i8_d2 (.clk(clk), .input_share0(d1_i8_s0), .input_share1(d1_i8_s1), .output_share0(d2_i8_s0), .output_share1(d2_i8_s1));
  reg_module u_reg_i9_d2 (.clk(clk), .input_share0(d1_i9_s0), .input_share1(d1_i9_s1), .output_share0(d2_i9_s0), .output_share1(d2_i9_s1));
  reg_module u_reg_t0_10_d2 (.clk(clk), .input_share0(d1_t0_10_s0), .input_share1(d1_t0_10_s1), .output_share0(d2_t0_10_s0), .output_share1(d2_t0_10_s1));
  reg_module u_reg_t0_11_d2 (.clk(clk), .input_share0(d1_t0_11_s0), .input_share1(d1_t0_11_s1), .output_share0(d2_t0_11_s0), .output_share1(d2_t0_11_s1));
  reg_module u_reg_t0_12_d2 (.clk(clk), .input_share0(d1_t0_12_s0), .input_share1(d1_t0_12_s1), .output_share0(d2_t0_12_s0), .output_share1(d2_t0_12_s1));
  reg_module u_reg_t0_13_d2 (.clk(clk), .input_share0(d1_t0_13_s0), .input_share1(d1_t0_13_s1), .output_share0(d2_t0_13_s0), .output_share1(d2_t0_13_s1));
  reg_module u_reg_t0_14_d2 (.clk(clk), .input_share0(d1_t0_14_s0), .input_share1(d1_t0_14_s1), .output_share0(d2_t0_14_s0), .output_share1(d2_t0_14_s1));
  reg_module u_reg_t0_15_d2 (.clk(clk), .input_share0(d1_t0_15_s0), .input_share1(d1_t0_15_s1), .output_share0(d2_t0_15_s0), .output_share1(d2_t0_15_s1));
  reg_module u_reg_t0_16_d2 (.clk(clk), .input_share0(d1_t0_16_s0), .input_share1(d1_t0_16_s1), .output_share0(d2_t0_16_s0), .output_share1(d2_t0_16_s1));
  reg_module u_reg_t0_17_d2 (.clk(clk), .input_share0(d1_t0_17_s0), .input_share1(d1_t0_17_s1), .output_share0(d2_t0_17_s0), .output_share1(d2_t0_17_s1));
  reg_module u_reg_t0_18_d2 (.clk(clk), .input_share0(d1_t0_18_s0), .input_share1(d1_t0_18_s1), .output_share0(d2_t0_18_s0), .output_share1(d2_t0_18_s1));
  reg_module u_reg_t0_19_d2 (.clk(clk), .input_share0(d1_t0_19_s0), .input_share1(d1_t0_19_s1), .output_share0(d2_t0_19_s0), .output_share1(d2_t0_19_s1));
  reg_module u_reg_t0_2_d2 (.clk(clk), .input_share0(d1_t0_2_s0), .input_share1(d1_t0_2_s1), .output_share0(d2_t0_2_s0), .output_share1(d2_t0_2_s1));
  reg_module u_reg_t0_20_d2 (.clk(clk), .input_share0(d1_t0_20_s0), .input_share1(d1_t0_20_s1), .output_share0(d2_t0_20_s0), .output_share1(d2_t0_20_s1));
  reg_module u_reg_t0_21_d2 (.clk(clk), .input_share0(d1_t0_21_s0), .input_share1(d1_t0_21_s1), .output_share0(d2_t0_21_s0), .output_share1(d2_t0_21_s1));
  reg_module u_reg_t0_22_d2 (.clk(clk), .input_share0(d1_t0_22_s0), .input_share1(d1_t0_22_s1), .output_share0(d2_t0_22_s0), .output_share1(d2_t0_22_s1));
  reg_module u_reg_t0_23_d2 (.clk(clk), .input_share0(d1_t0_23_s0), .input_share1(d1_t0_23_s1), .output_share0(d2_t0_23_s0), .output_share1(d2_t0_23_s1));
  reg_module u_reg_t0_24_d2 (.clk(clk), .input_share0(d1_t0_24_s0), .input_share1(d1_t0_24_s1), .output_share0(d2_t0_24_s0), .output_share1(d2_t0_24_s1));
  reg_module u_reg_t0_25_d2 (.clk(clk), .input_share0(d1_t0_25_s0), .input_share1(d1_t0_25_s1), .output_share0(d2_t0_25_s0), .output_share1(d2_t0_25_s1));
  reg_module u_reg_t0_26_d2 (.clk(clk), .input_share0(d1_t0_26_s0), .input_share1(d1_t0_26_s1), .output_share0(d2_t0_26_s0), .output_share1(d2_t0_26_s1));
  reg_module u_reg_t0_27_d2 (.clk(clk), .input_share0(d1_t0_27_s0), .input_share1(d1_t0_27_s1), .output_share0(d2_t0_27_s0), .output_share1(d2_t0_27_s1));
  reg_module u_reg_t0_28_d2 (.clk(clk), .input_share0(d1_t0_28_s0), .input_share1(d1_t0_28_s1), .output_share0(d2_t0_28_s0), .output_share1(d2_t0_28_s1));
  reg_module u_reg_t0_29_d2 (.clk(clk), .input_share0(d1_t0_29_s0), .input_share1(d1_t0_29_s1), .output_share0(d2_t0_29_s0), .output_share1(d2_t0_29_s1));
  reg_module u_reg_t0_3_d2 (.clk(clk), .input_share0(d1_t0_3_s0), .input_share1(d1_t0_3_s1), .output_share0(d2_t0_3_s0), .output_share1(d2_t0_3_s1));
  reg_module u_reg_t0_30_d2 (.clk(clk), .input_share0(d1_t0_30_s0), .input_share1(d1_t0_30_s1), .output_share0(d2_t0_30_s0), .output_share1(d2_t0_30_s1));
  reg_module u_reg_t0_31_d2 (.clk(clk), .input_share0(d1_t0_31_s0), .input_share1(d1_t0_31_s1), .output_share0(d2_t0_31_s0), .output_share1(d2_t0_31_s1));
  reg_module u_reg_t0_4_d2 (.clk(clk), .input_share0(d1_t0_4_s0), .input_share1(d1_t0_4_s1), .output_share0(d2_t0_4_s0), .output_share1(d2_t0_4_s1));
  reg_module u_reg_t0_5_d2 (.clk(clk), .input_share0(d1_t0_5_s0), .input_share1(d1_t0_5_s1), .output_share0(d2_t0_5_s0), .output_share1(d2_t0_5_s1));
  reg_module u_reg_t0_6_d2 (.clk(clk), .input_share0(d1_t0_6_s0), .input_share1(d1_t0_6_s1), .output_share0(d2_t0_6_s0), .output_share1(d2_t0_6_s1));
  reg_module u_reg_t0_7_d2 (.clk(clk), .input_share0(d1_t0_7_s0), .input_share1(d1_t0_7_s1), .output_share0(d2_t0_7_s0), .output_share1(d2_t0_7_s1));
  reg_module u_reg_t0_8_d2 (.clk(clk), .input_share0(d1_t0_8_s0), .input_share1(d1_t0_8_s1), .output_share0(d2_t0_8_s0), .output_share1(d2_t0_8_s1));
  reg_module u_reg_t0_9_d2 (.clk(clk), .input_share0(d1_t0_9_s0), .input_share1(d1_t0_9_s1), .output_share0(d2_t0_9_s0), .output_share1(d2_t0_9_s1));
  xor_module u_xor_c2_d2 (.x_share0(d2_i1_s0), .x_share1(d2_i1_s1), .y_share0(d2_t2_1_s0), .y_share1(d2_t2_1_s1), .z_share0(d2_c2_s0), .z_share1(d2_c2_s1));
  xor_module u_xor_o2_d2 (.x_share0(d2_t0_2_s0), .x_share1(d2_t0_2_s1), .y_share0(d2_c2_s0), .y_share1(d2_c2_s1), .z_share0(d2_o2_s0), .z_share1(d2_o2_s1));
  xor_module u_xor_t1_2_d2 (.x_share0(d2_i2_s0), .x_share1(d2_i2_s1), .y_share0(d2_c2_s0), .y_share1(d2_c2_s1), .z_share0(d2_t1_2_s0), .z_share1(d2_t1_2_s1));
  and_module u_and_t2_1_d2 (.clk(clk), .x_share0(d1_t0_1_s0), .x_share1(d1_t0_1_s1), .y_share0(d1_t1_1_s0), .y_share1(d1_t1_1_s1), .rand(r_t2_1), .z_share0(d2_t2_1_s0), .z_share1(d2_t2_1_s1));
  assign r_t2_1 = stage2_share0[2];
  reg_module u_reg_i10_d3 (.clk(clk), .input_share0(d2_i10_s0), .input_share1(d2_i10_s1), .output_share0(d3_i10_s0), .output_share1(d3_i10_s1));
  reg_module u_reg_i11_d3 (.clk(clk), .input_share0(d2_i11_s0), .input_share1(d2_i11_s1), .output_share0(d3_i11_s0), .output_share1(d3_i11_s1));
  reg_module u_reg_i12_d3 (.clk(clk), .input_share0(d2_i12_s0), .input_share1(d2_i12_s1), .output_share0(d3_i12_s0), .output_share1(d3_i12_s1));
  reg_module u_reg_i13_d3 (.clk(clk), .input_share0(d2_i13_s0), .input_share1(d2_i13_s1), .output_share0(d3_i13_s0), .output_share1(d3_i13_s1));
  reg_module u_reg_i14_d3 (.clk(clk), .input_share0(d2_i14_s0), .input_share1(d2_i14_s1), .output_share0(d3_i14_s0), .output_share1(d3_i14_s1));
  reg_module u_reg_i15_d3 (.clk(clk), .input_share0(d2_i15_s0), .input_share1(d2_i15_s1), .output_share0(d3_i15_s0), .output_share1(d3_i15_s1));
  reg_module u_reg_i16_d3 (.clk(clk), .input_share0(d2_i16_s0), .input_share1(d2_i16_s1), .output_share0(d3_i16_s0), .output_share1(d3_i16_s1));
  reg_module u_reg_i17_d3 (.clk(clk), .input_share0(d2_i17_s0), .input_share1(d2_i17_s1), .output_share0(d3_i17_s0), .output_share1(d3_i17_s1));
  reg_module u_reg_i18_d3 (.clk(clk), .input_share0(d2_i18_s0), .input_share1(d2_i18_s1), .output_share0(d3_i18_s0), .output_share1(d3_i18_s1));
  reg_module u_reg_i19_d3 (.clk(clk), .input_share0(d2_i19_s0), .input_share1(d2_i19_s1), .output_share0(d3_i19_s0), .output_share1(d3_i19_s1));
  reg_module u_reg_i2_d3 (.clk(clk), .input_share0(d2_i2_s0), .input_share1(d2_i2_s1), .output_share0(d3_i2_s0), .output_share1(d3_i2_s1));
  reg_module u_reg_i20_d3 (.clk(clk), .input_share0(d2_i20_s0), .input_share1(d2_i20_s1), .output_share0(d3_i20_s0), .output_share1(d3_i20_s1));
  reg_module u_reg_i21_d3 (.clk(clk), .input_share0(d2_i21_s0), .input_share1(d2_i21_s1), .output_share0(d3_i21_s0), .output_share1(d3_i21_s1));
  reg_module u_reg_i22_d3 (.clk(clk), .input_share0(d2_i22_s0), .input_share1(d2_i22_s1), .output_share0(d3_i22_s0), .output_share1(d3_i22_s1));
  reg_module u_reg_i23_d3 (.clk(clk), .input_share0(d2_i23_s0), .input_share1(d2_i23_s1), .output_share0(d3_i23_s0), .output_share1(d3_i23_s1));
  reg_module u_reg_i24_d3 (.clk(clk), .input_share0(d2_i24_s0), .input_share1(d2_i24_s1), .output_share0(d3_i24_s0), .output_share1(d3_i24_s1));
  reg_module u_reg_i25_d3 (.clk(clk), .input_share0(d2_i25_s0), .input_share1(d2_i25_s1), .output_share0(d3_i25_s0), .output_share1(d3_i25_s1));
  reg_module u_reg_i26_d3 (.clk(clk), .input_share0(d2_i26_s0), .input_share1(d2_i26_s1), .output_share0(d3_i26_s0), .output_share1(d3_i26_s1));
  reg_module u_reg_i27_d3 (.clk(clk), .input_share0(d2_i27_s0), .input_share1(d2_i27_s1), .output_share0(d3_i27_s0), .output_share1(d3_i27_s1));
  reg_module u_reg_i28_d3 (.clk(clk), .input_share0(d2_i28_s0), .input_share1(d2_i28_s1), .output_share0(d3_i28_s0), .output_share1(d3_i28_s1));
  reg_module u_reg_i29_d3 (.clk(clk), .input_share0(d2_i29_s0), .input_share1(d2_i29_s1), .output_share0(d3_i29_s0), .output_share1(d3_i29_s1));
  reg_module u_reg_i3_d3 (.clk(clk), .input_share0(d2_i3_s0), .input_share1(d2_i3_s1), .output_share0(d3_i3_s0), .output_share1(d3_i3_s1));
  reg_module u_reg_i30_d3 (.clk(clk), .input_share0(d2_i30_s0), .input_share1(d2_i30_s1), .output_share0(d3_i30_s0), .output_share1(d3_i30_s1));
  reg_module u_reg_i4_d3 (.clk(clk), .input_share0(d2_i4_s0), .input_share1(d2_i4_s1), .output_share0(d3_i4_s0), .output_share1(d3_i4_s1));
  reg_module u_reg_i5_d3 (.clk(clk), .input_share0(d2_i5_s0), .input_share1(d2_i5_s1), .output_share0(d3_i5_s0), .output_share1(d3_i5_s1));
  reg_module u_reg_i6_d3 (.clk(clk), .input_share0(d2_i6_s0), .input_share1(d2_i6_s1), .output_share0(d3_i6_s0), .output_share1(d3_i6_s1));
  reg_module u_reg_i7_d3 (.clk(clk), .input_share0(d2_i7_s0), .input_share1(d2_i7_s1), .output_share0(d3_i7_s0), .output_share1(d3_i7_s1));
  reg_module u_reg_i8_d3 (.clk(clk), .input_share0(d2_i8_s0), .input_share1(d2_i8_s1), .output_share0(d3_i8_s0), .output_share1(d3_i8_s1));
  reg_module u_reg_i9_d3 (.clk(clk), .input_share0(d2_i9_s0), .input_share1(d2_i9_s1), .output_share0(d3_i9_s0), .output_share1(d3_i9_s1));
  reg_module u_reg_t0_10_d3 (.clk(clk), .input_share0(d2_t0_10_s0), .input_share1(d2_t0_10_s1), .output_share0(d3_t0_10_s0), .output_share1(d3_t0_10_s1));
  reg_module u_reg_t0_11_d3 (.clk(clk), .input_share0(d2_t0_11_s0), .input_share1(d2_t0_11_s1), .output_share0(d3_t0_11_s0), .output_share1(d3_t0_11_s1));
  reg_module u_reg_t0_12_d3 (.clk(clk), .input_share0(d2_t0_12_s0), .input_share1(d2_t0_12_s1), .output_share0(d3_t0_12_s0), .output_share1(d3_t0_12_s1));
  reg_module u_reg_t0_13_d3 (.clk(clk), .input_share0(d2_t0_13_s0), .input_share1(d2_t0_13_s1), .output_share0(d3_t0_13_s0), .output_share1(d3_t0_13_s1));
  reg_module u_reg_t0_14_d3 (.clk(clk), .input_share0(d2_t0_14_s0), .input_share1(d2_t0_14_s1), .output_share0(d3_t0_14_s0), .output_share1(d3_t0_14_s1));
  reg_module u_reg_t0_15_d3 (.clk(clk), .input_share0(d2_t0_15_s0), .input_share1(d2_t0_15_s1), .output_share0(d3_t0_15_s0), .output_share1(d3_t0_15_s1));
  reg_module u_reg_t0_16_d3 (.clk(clk), .input_share0(d2_t0_16_s0), .input_share1(d2_t0_16_s1), .output_share0(d3_t0_16_s0), .output_share1(d3_t0_16_s1));
  reg_module u_reg_t0_17_d3 (.clk(clk), .input_share0(d2_t0_17_s0), .input_share1(d2_t0_17_s1), .output_share0(d3_t0_17_s0), .output_share1(d3_t0_17_s1));
  reg_module u_reg_t0_18_d3 (.clk(clk), .input_share0(d2_t0_18_s0), .input_share1(d2_t0_18_s1), .output_share0(d3_t0_18_s0), .output_share1(d3_t0_18_s1));
  reg_module u_reg_t0_19_d3 (.clk(clk), .input_share0(d2_t0_19_s0), .input_share1(d2_t0_19_s1), .output_share0(d3_t0_19_s0), .output_share1(d3_t0_19_s1));
  reg_module u_reg_t0_20_d3 (.clk(clk), .input_share0(d2_t0_20_s0), .input_share1(d2_t0_20_s1), .output_share0(d3_t0_20_s0), .output_share1(d3_t0_20_s1));
  reg_module u_reg_t0_21_d3 (.clk(clk), .input_share0(d2_t0_21_s0), .input_share1(d2_t0_21_s1), .output_share0(d3_t0_21_s0), .output_share1(d3_t0_21_s1));
  reg_module u_reg_t0_22_d3 (.clk(clk), .input_share0(d2_t0_22_s0), .input_share1(d2_t0_22_s1), .output_share0(d3_t0_22_s0), .output_share1(d3_t0_22_s1));
  reg_module u_reg_t0_23_d3 (.clk(clk), .input_share0(d2_t0_23_s0), .input_share1(d2_t0_23_s1), .output_share0(d3_t0_23_s0), .output_share1(d3_t0_23_s1));
  reg_module u_reg_t0_24_d3 (.clk(clk), .input_share0(d2_t0_24_s0), .input_share1(d2_t0_24_s1), .output_share0(d3_t0_24_s0), .output_share1(d3_t0_24_s1));
  reg_module u_reg_t0_25_d3 (.clk(clk), .input_share0(d2_t0_25_s0), .input_share1(d2_t0_25_s1), .output_share0(d3_t0_25_s0), .output_share1(d3_t0_25_s1));
  reg_module u_reg_t0_26_d3 (.clk(clk), .input_share0(d2_t0_26_s0), .input_share1(d2_t0_26_s1), .output_share0(d3_t0_26_s0), .output_share1(d3_t0_26_s1));
  reg_module u_reg_t0_27_d3 (.clk(clk), .input_share0(d2_t0_27_s0), .input_share1(d2_t0_27_s1), .output_share0(d3_t0_27_s0), .output_share1(d3_t0_27_s1));
  reg_module u_reg_t0_28_d3 (.clk(clk), .input_share0(d2_t0_28_s0), .input_share1(d2_t0_28_s1), .output_share0(d3_t0_28_s0), .output_share1(d3_t0_28_s1));
  reg_module u_reg_t0_29_d3 (.clk(clk), .input_share0(d2_t0_29_s0), .input_share1(d2_t0_29_s1), .output_share0(d3_t0_29_s0), .output_share1(d3_t0_29_s1));
  reg_module u_reg_t0_3_d3 (.clk(clk), .input_share0(d2_t0_3_s0), .input_share1(d2_t0_3_s1), .output_share0(d3_t0_3_s0), .output_share1(d3_t0_3_s1));
  reg_module u_reg_t0_30_d3 (.clk(clk), .input_share0(d2_t0_30_s0), .input_share1(d2_t0_30_s1), .output_share0(d3_t0_30_s0), .output_share1(d3_t0_30_s1));
  reg_module u_reg_t0_31_d3 (.clk(clk), .input_share0(d2_t0_31_s0), .input_share1(d2_t0_31_s1), .output_share0(d3_t0_31_s0), .output_share1(d3_t0_31_s1));
  reg_module u_reg_t0_4_d3 (.clk(clk), .input_share0(d2_t0_4_s0), .input_share1(d2_t0_4_s1), .output_share0(d3_t0_4_s0), .output_share1(d3_t0_4_s1));
  reg_module u_reg_t0_5_d3 (.clk(clk), .input_share0(d2_t0_5_s0), .input_share1(d2_t0_5_s1), .output_share0(d3_t0_5_s0), .output_share1(d3_t0_5_s1));
  reg_module u_reg_t0_6_d3 (.clk(clk), .input_share0(d2_t0_6_s0), .input_share1(d2_t0_6_s1), .output_share0(d3_t0_6_s0), .output_share1(d3_t0_6_s1));
  reg_module u_reg_t0_7_d3 (.clk(clk), .input_share0(d2_t0_7_s0), .input_share1(d2_t0_7_s1), .output_share0(d3_t0_7_s0), .output_share1(d3_t0_7_s1));
  reg_module u_reg_t0_8_d3 (.clk(clk), .input_share0(d2_t0_8_s0), .input_share1(d2_t0_8_s1), .output_share0(d3_t0_8_s0), .output_share1(d3_t0_8_s1));
  reg_module u_reg_t0_9_d3 (.clk(clk), .input_share0(d2_t0_9_s0), .input_share1(d2_t0_9_s1), .output_share0(d3_t0_9_s0), .output_share1(d3_t0_9_s1));
  xor_module u_xor_c3_d3 (.x_share0(d3_i2_s0), .x_share1(d3_i2_s1), .y_share0(d3_t2_2_s0), .y_share1(d3_t2_2_s1), .z_share0(d3_c3_s0), .z_share1(d3_c3_s1));
  xor_module u_xor_o3_d3 (.x_share0(d3_t0_3_s0), .x_share1(d3_t0_3_s1), .y_share0(d3_c3_s0), .y_share1(d3_c3_s1), .z_share0(d3_o3_s0), .z_share1(d3_o3_s1));
  xor_module u_xor_t1_3_d3 (.x_share0(d3_i3_s0), .x_share1(d3_i3_s1), .y_share0(d3_c3_s0), .y_share1(d3_c3_s1), .z_share0(d3_t1_3_s0), .z_share1(d3_t1_3_s1));
  and_module u_and_t2_2_d3 (.clk(clk), .x_share0(d2_t0_2_s0), .x_share1(d2_t0_2_s1), .y_share0(d2_t1_2_s0), .y_share1(d2_t1_2_s1), .rand(r_t2_2), .z_share0(d3_t2_2_s0), .z_share1(d3_t2_2_s1));
  assign r_t2_2 = stage3_share0[0];
  reg_module u_reg_i10_d4 (.clk(clk), .input_share0(d3_i10_s0), .input_share1(d3_i10_s1), .output_share0(d4_i10_s0), .output_share1(d4_i10_s1));
  reg_module u_reg_i11_d4 (.clk(clk), .input_share0(d3_i11_s0), .input_share1(d3_i11_s1), .output_share0(d4_i11_s0), .output_share1(d4_i11_s1));
  reg_module u_reg_i12_d4 (.clk(clk), .input_share0(d3_i12_s0), .input_share1(d3_i12_s1), .output_share0(d4_i12_s0), .output_share1(d4_i12_s1));
  reg_module u_reg_i13_d4 (.clk(clk), .input_share0(d3_i13_s0), .input_share1(d3_i13_s1), .output_share0(d4_i13_s0), .output_share1(d4_i13_s1));
  reg_module u_reg_i14_d4 (.clk(clk), .input_share0(d3_i14_s0), .input_share1(d3_i14_s1), .output_share0(d4_i14_s0), .output_share1(d4_i14_s1));
  reg_module u_reg_i15_d4 (.clk(clk), .input_share0(d3_i15_s0), .input_share1(d3_i15_s1), .output_share0(d4_i15_s0), .output_share1(d4_i15_s1));
  reg_module u_reg_i16_d4 (.clk(clk), .input_share0(d3_i16_s0), .input_share1(d3_i16_s1), .output_share0(d4_i16_s0), .output_share1(d4_i16_s1));
  reg_module u_reg_i17_d4 (.clk(clk), .input_share0(d3_i17_s0), .input_share1(d3_i17_s1), .output_share0(d4_i17_s0), .output_share1(d4_i17_s1));
  reg_module u_reg_i18_d4 (.clk(clk), .input_share0(d3_i18_s0), .input_share1(d3_i18_s1), .output_share0(d4_i18_s0), .output_share1(d4_i18_s1));
  reg_module u_reg_i19_d4 (.clk(clk), .input_share0(d3_i19_s0), .input_share1(d3_i19_s1), .output_share0(d4_i19_s0), .output_share1(d4_i19_s1));
  reg_module u_reg_i20_d4 (.clk(clk), .input_share0(d3_i20_s0), .input_share1(d3_i20_s1), .output_share0(d4_i20_s0), .output_share1(d4_i20_s1));
  reg_module u_reg_i21_d4 (.clk(clk), .input_share0(d3_i21_s0), .input_share1(d3_i21_s1), .output_share0(d4_i21_s0), .output_share1(d4_i21_s1));
  reg_module u_reg_i22_d4 (.clk(clk), .input_share0(d3_i22_s0), .input_share1(d3_i22_s1), .output_share0(d4_i22_s0), .output_share1(d4_i22_s1));
  reg_module u_reg_i23_d4 (.clk(clk), .input_share0(d3_i23_s0), .input_share1(d3_i23_s1), .output_share0(d4_i23_s0), .output_share1(d4_i23_s1));
  reg_module u_reg_i24_d4 (.clk(clk), .input_share0(d3_i24_s0), .input_share1(d3_i24_s1), .output_share0(d4_i24_s0), .output_share1(d4_i24_s1));
  reg_module u_reg_i25_d4 (.clk(clk), .input_share0(d3_i25_s0), .input_share1(d3_i25_s1), .output_share0(d4_i25_s0), .output_share1(d4_i25_s1));
  reg_module u_reg_i26_d4 (.clk(clk), .input_share0(d3_i26_s0), .input_share1(d3_i26_s1), .output_share0(d4_i26_s0), .output_share1(d4_i26_s1));
  reg_module u_reg_i27_d4 (.clk(clk), .input_share0(d3_i27_s0), .input_share1(d3_i27_s1), .output_share0(d4_i27_s0), .output_share1(d4_i27_s1));
  reg_module u_reg_i28_d4 (.clk(clk), .input_share0(d3_i28_s0), .input_share1(d3_i28_s1), .output_share0(d4_i28_s0), .output_share1(d4_i28_s1));
  reg_module u_reg_i29_d4 (.clk(clk), .input_share0(d3_i29_s0), .input_share1(d3_i29_s1), .output_share0(d4_i29_s0), .output_share1(d4_i29_s1));
  reg_module u_reg_i3_d4 (.clk(clk), .input_share0(d3_i3_s0), .input_share1(d3_i3_s1), .output_share0(d4_i3_s0), .output_share1(d4_i3_s1));
  reg_module u_reg_i30_d4 (.clk(clk), .input_share0(d3_i30_s0), .input_share1(d3_i30_s1), .output_share0(d4_i30_s0), .output_share1(d4_i30_s1));
  reg_module u_reg_i4_d4 (.clk(clk), .input_share0(d3_i4_s0), .input_share1(d3_i4_s1), .output_share0(d4_i4_s0), .output_share1(d4_i4_s1));
  reg_module u_reg_i5_d4 (.clk(clk), .input_share0(d3_i5_s0), .input_share1(d3_i5_s1), .output_share0(d4_i5_s0), .output_share1(d4_i5_s1));
  reg_module u_reg_i6_d4 (.clk(clk), .input_share0(d3_i6_s0), .input_share1(d3_i6_s1), .output_share0(d4_i6_s0), .output_share1(d4_i6_s1));
  reg_module u_reg_i7_d4 (.clk(clk), .input_share0(d3_i7_s0), .input_share1(d3_i7_s1), .output_share0(d4_i7_s0), .output_share1(d4_i7_s1));
  reg_module u_reg_i8_d4 (.clk(clk), .input_share0(d3_i8_s0), .input_share1(d3_i8_s1), .output_share0(d4_i8_s0), .output_share1(d4_i8_s1));
  reg_module u_reg_i9_d4 (.clk(clk), .input_share0(d3_i9_s0), .input_share1(d3_i9_s1), .output_share0(d4_i9_s0), .output_share1(d4_i9_s1));
  reg_module u_reg_t0_10_d4 (.clk(clk), .input_share0(d3_t0_10_s0), .input_share1(d3_t0_10_s1), .output_share0(d4_t0_10_s0), .output_share1(d4_t0_10_s1));
  reg_module u_reg_t0_11_d4 (.clk(clk), .input_share0(d3_t0_11_s0), .input_share1(d3_t0_11_s1), .output_share0(d4_t0_11_s0), .output_share1(d4_t0_11_s1));
  reg_module u_reg_t0_12_d4 (.clk(clk), .input_share0(d3_t0_12_s0), .input_share1(d3_t0_12_s1), .output_share0(d4_t0_12_s0), .output_share1(d4_t0_12_s1));
  reg_module u_reg_t0_13_d4 (.clk(clk), .input_share0(d3_t0_13_s0), .input_share1(d3_t0_13_s1), .output_share0(d4_t0_13_s0), .output_share1(d4_t0_13_s1));
  reg_module u_reg_t0_14_d4 (.clk(clk), .input_share0(d3_t0_14_s0), .input_share1(d3_t0_14_s1), .output_share0(d4_t0_14_s0), .output_share1(d4_t0_14_s1));
  reg_module u_reg_t0_15_d4 (.clk(clk), .input_share0(d3_t0_15_s0), .input_share1(d3_t0_15_s1), .output_share0(d4_t0_15_s0), .output_share1(d4_t0_15_s1));
  reg_module u_reg_t0_16_d4 (.clk(clk), .input_share0(d3_t0_16_s0), .input_share1(d3_t0_16_s1), .output_share0(d4_t0_16_s0), .output_share1(d4_t0_16_s1));
  reg_module u_reg_t0_17_d4 (.clk(clk), .input_share0(d3_t0_17_s0), .input_share1(d3_t0_17_s1), .output_share0(d4_t0_17_s0), .output_share1(d4_t0_17_s1));
  reg_module u_reg_t0_18_d4 (.clk(clk), .input_share0(d3_t0_18_s0), .input_share1(d3_t0_18_s1), .output_share0(d4_t0_18_s0), .output_share1(d4_t0_18_s1));
  reg_module u_reg_t0_19_d4 (.clk(clk), .input_share0(d3_t0_19_s0), .input_share1(d3_t0_19_s1), .output_share0(d4_t0_19_s0), .output_share1(d4_t0_19_s1));
  reg_module u_reg_t0_20_d4 (.clk(clk), .input_share0(d3_t0_20_s0), .input_share1(d3_t0_20_s1), .output_share0(d4_t0_20_s0), .output_share1(d4_t0_20_s1));
  reg_module u_reg_t0_21_d4 (.clk(clk), .input_share0(d3_t0_21_s0), .input_share1(d3_t0_21_s1), .output_share0(d4_t0_21_s0), .output_share1(d4_t0_21_s1));
  reg_module u_reg_t0_22_d4 (.clk(clk), .input_share0(d3_t0_22_s0), .input_share1(d3_t0_22_s1), .output_share0(d4_t0_22_s0), .output_share1(d4_t0_22_s1));
  reg_module u_reg_t0_23_d4 (.clk(clk), .input_share0(d3_t0_23_s0), .input_share1(d3_t0_23_s1), .output_share0(d4_t0_23_s0), .output_share1(d4_t0_23_s1));
  reg_module u_reg_t0_24_d4 (.clk(clk), .input_share0(d3_t0_24_s0), .input_share1(d3_t0_24_s1), .output_share0(d4_t0_24_s0), .output_share1(d4_t0_24_s1));
  reg_module u_reg_t0_25_d4 (.clk(clk), .input_share0(d3_t0_25_s0), .input_share1(d3_t0_25_s1), .output_share0(d4_t0_25_s0), .output_share1(d4_t0_25_s1));
  reg_module u_reg_t0_26_d4 (.clk(clk), .input_share0(d3_t0_26_s0), .input_share1(d3_t0_26_s1), .output_share0(d4_t0_26_s0), .output_share1(d4_t0_26_s1));
  reg_module u_reg_t0_27_d4 (.clk(clk), .input_share0(d3_t0_27_s0), .input_share1(d3_t0_27_s1), .output_share0(d4_t0_27_s0), .output_share1(d4_t0_27_s1));
  reg_module u_reg_t0_28_d4 (.clk(clk), .input_share0(d3_t0_28_s0), .input_share1(d3_t0_28_s1), .output_share0(d4_t0_28_s0), .output_share1(d4_t0_28_s1));
  reg_module u_reg_t0_29_d4 (.clk(clk), .input_share0(d3_t0_29_s0), .input_share1(d3_t0_29_s1), .output_share0(d4_t0_29_s0), .output_share1(d4_t0_29_s1));
  reg_module u_reg_t0_30_d4 (.clk(clk), .input_share0(d3_t0_30_s0), .input_share1(d3_t0_30_s1), .output_share0(d4_t0_30_s0), .output_share1(d4_t0_30_s1));
  reg_module u_reg_t0_31_d4 (.clk(clk), .input_share0(d3_t0_31_s0), .input_share1(d3_t0_31_s1), .output_share0(d4_t0_31_s0), .output_share1(d4_t0_31_s1));
  reg_module u_reg_t0_4_d4 (.clk(clk), .input_share0(d3_t0_4_s0), .input_share1(d3_t0_4_s1), .output_share0(d4_t0_4_s0), .output_share1(d4_t0_4_s1));
  reg_module u_reg_t0_5_d4 (.clk(clk), .input_share0(d3_t0_5_s0), .input_share1(d3_t0_5_s1), .output_share0(d4_t0_5_s0), .output_share1(d4_t0_5_s1));
  reg_module u_reg_t0_6_d4 (.clk(clk), .input_share0(d3_t0_6_s0), .input_share1(d3_t0_6_s1), .output_share0(d4_t0_6_s0), .output_share1(d4_t0_6_s1));
  reg_module u_reg_t0_7_d4 (.clk(clk), .input_share0(d3_t0_7_s0), .input_share1(d3_t0_7_s1), .output_share0(d4_t0_7_s0), .output_share1(d4_t0_7_s1));
  reg_module u_reg_t0_8_d4 (.clk(clk), .input_share0(d3_t0_8_s0), .input_share1(d3_t0_8_s1), .output_share0(d4_t0_8_s0), .output_share1(d4_t0_8_s1));
  reg_module u_reg_t0_9_d4 (.clk(clk), .input_share0(d3_t0_9_s0), .input_share1(d3_t0_9_s1), .output_share0(d4_t0_9_s0), .output_share1(d4_t0_9_s1));
  xor_module u_xor_c4_d4 (.x_share0(d4_i3_s0), .x_share1(d4_i3_s1), .y_share0(d4_t2_3_s0), .y_share1(d4_t2_3_s1), .z_share0(d4_c4_s0), .z_share1(d4_c4_s1));
  xor_module u_xor_o4_d4 (.x_share0(d4_t0_4_s0), .x_share1(d4_t0_4_s1), .y_share0(d4_c4_s0), .y_share1(d4_c4_s1), .z_share0(d4_o4_s0), .z_share1(d4_o4_s1));
  xor_module u_xor_t1_4_d4 (.x_share0(d4_i4_s0), .x_share1(d4_i4_s1), .y_share0(d4_c4_s0), .y_share1(d4_c4_s1), .z_share0(d4_t1_4_s0), .z_share1(d4_t1_4_s1));
  and_module u_and_t2_3_d4 (.clk(clk), .x_share0(d3_t0_3_s0), .x_share1(d3_t0_3_s1), .y_share0(d3_t1_3_s0), .y_share1(d3_t1_3_s1), .rand(r_t2_3), .z_share0(d4_t2_3_s0), .z_share1(d4_t2_3_s1));
  assign r_t2_3 = stage4_share0[1];
  reg_module u_reg_i10_d5 (.clk(clk), .input_share0(d4_i10_s0), .input_share1(d4_i10_s1), .output_share0(d5_i10_s0), .output_share1(d5_i10_s1));
  reg_module u_reg_i11_d5 (.clk(clk), .input_share0(d4_i11_s0), .input_share1(d4_i11_s1), .output_share0(d5_i11_s0), .output_share1(d5_i11_s1));
  reg_module u_reg_i12_d5 (.clk(clk), .input_share0(d4_i12_s0), .input_share1(d4_i12_s1), .output_share0(d5_i12_s0), .output_share1(d5_i12_s1));
  reg_module u_reg_i13_d5 (.clk(clk), .input_share0(d4_i13_s0), .input_share1(d4_i13_s1), .output_share0(d5_i13_s0), .output_share1(d5_i13_s1));
  reg_module u_reg_i14_d5 (.clk(clk), .input_share0(d4_i14_s0), .input_share1(d4_i14_s1), .output_share0(d5_i14_s0), .output_share1(d5_i14_s1));
  reg_module u_reg_i15_d5 (.clk(clk), .input_share0(d4_i15_s0), .input_share1(d4_i15_s1), .output_share0(d5_i15_s0), .output_share1(d5_i15_s1));
  reg_module u_reg_i16_d5 (.clk(clk), .input_share0(d4_i16_s0), .input_share1(d4_i16_s1), .output_share0(d5_i16_s0), .output_share1(d5_i16_s1));
  reg_module u_reg_i17_d5 (.clk(clk), .input_share0(d4_i17_s0), .input_share1(d4_i17_s1), .output_share0(d5_i17_s0), .output_share1(d5_i17_s1));
  reg_module u_reg_i18_d5 (.clk(clk), .input_share0(d4_i18_s0), .input_share1(d4_i18_s1), .output_share0(d5_i18_s0), .output_share1(d5_i18_s1));
  reg_module u_reg_i19_d5 (.clk(clk), .input_share0(d4_i19_s0), .input_share1(d4_i19_s1), .output_share0(d5_i19_s0), .output_share1(d5_i19_s1));
  reg_module u_reg_i20_d5 (.clk(clk), .input_share0(d4_i20_s0), .input_share1(d4_i20_s1), .output_share0(d5_i20_s0), .output_share1(d5_i20_s1));
  reg_module u_reg_i21_d5 (.clk(clk), .input_share0(d4_i21_s0), .input_share1(d4_i21_s1), .output_share0(d5_i21_s0), .output_share1(d5_i21_s1));
  reg_module u_reg_i22_d5 (.clk(clk), .input_share0(d4_i22_s0), .input_share1(d4_i22_s1), .output_share0(d5_i22_s0), .output_share1(d5_i22_s1));
  reg_module u_reg_i23_d5 (.clk(clk), .input_share0(d4_i23_s0), .input_share1(d4_i23_s1), .output_share0(d5_i23_s0), .output_share1(d5_i23_s1));
  reg_module u_reg_i24_d5 (.clk(clk), .input_share0(d4_i24_s0), .input_share1(d4_i24_s1), .output_share0(d5_i24_s0), .output_share1(d5_i24_s1));
  reg_module u_reg_i25_d5 (.clk(clk), .input_share0(d4_i25_s0), .input_share1(d4_i25_s1), .output_share0(d5_i25_s0), .output_share1(d5_i25_s1));
  reg_module u_reg_i26_d5 (.clk(clk), .input_share0(d4_i26_s0), .input_share1(d4_i26_s1), .output_share0(d5_i26_s0), .output_share1(d5_i26_s1));
  reg_module u_reg_i27_d5 (.clk(clk), .input_share0(d4_i27_s0), .input_share1(d4_i27_s1), .output_share0(d5_i27_s0), .output_share1(d5_i27_s1));
  reg_module u_reg_i28_d5 (.clk(clk), .input_share0(d4_i28_s0), .input_share1(d4_i28_s1), .output_share0(d5_i28_s0), .output_share1(d5_i28_s1));
  reg_module u_reg_i29_d5 (.clk(clk), .input_share0(d4_i29_s0), .input_share1(d4_i29_s1), .output_share0(d5_i29_s0), .output_share1(d5_i29_s1));
  reg_module u_reg_i30_d5 (.clk(clk), .input_share0(d4_i30_s0), .input_share1(d4_i30_s1), .output_share0(d5_i30_s0), .output_share1(d5_i30_s1));
  reg_module u_reg_i4_d5 (.clk(clk), .input_share0(d4_i4_s0), .input_share1(d4_i4_s1), .output_share0(d5_i4_s0), .output_share1(d5_i4_s1));
  reg_module u_reg_i5_d5 (.clk(clk), .input_share0(d4_i5_s0), .input_share1(d4_i5_s1), .output_share0(d5_i5_s0), .output_share1(d5_i5_s1));
  reg_module u_reg_i6_d5 (.clk(clk), .input_share0(d4_i6_s0), .input_share1(d4_i6_s1), .output_share0(d5_i6_s0), .output_share1(d5_i6_s1));
  reg_module u_reg_i7_d5 (.clk(clk), .input_share0(d4_i7_s0), .input_share1(d4_i7_s1), .output_share0(d5_i7_s0), .output_share1(d5_i7_s1));
  reg_module u_reg_i8_d5 (.clk(clk), .input_share0(d4_i8_s0), .input_share1(d4_i8_s1), .output_share0(d5_i8_s0), .output_share1(d5_i8_s1));
  reg_module u_reg_i9_d5 (.clk(clk), .input_share0(d4_i9_s0), .input_share1(d4_i9_s1), .output_share0(d5_i9_s0), .output_share1(d5_i9_s1));
  reg_module u_reg_t0_10_d5 (.clk(clk), .input_share0(d4_t0_10_s0), .input_share1(d4_t0_10_s1), .output_share0(d5_t0_10_s0), .output_share1(d5_t0_10_s1));
  reg_module u_reg_t0_11_d5 (.clk(clk), .input_share0(d4_t0_11_s0), .input_share1(d4_t0_11_s1), .output_share0(d5_t0_11_s0), .output_share1(d5_t0_11_s1));
  reg_module u_reg_t0_12_d5 (.clk(clk), .input_share0(d4_t0_12_s0), .input_share1(d4_t0_12_s1), .output_share0(d5_t0_12_s0), .output_share1(d5_t0_12_s1));
  reg_module u_reg_t0_13_d5 (.clk(clk), .input_share0(d4_t0_13_s0), .input_share1(d4_t0_13_s1), .output_share0(d5_t0_13_s0), .output_share1(d5_t0_13_s1));
  reg_module u_reg_t0_14_d5 (.clk(clk), .input_share0(d4_t0_14_s0), .input_share1(d4_t0_14_s1), .output_share0(d5_t0_14_s0), .output_share1(d5_t0_14_s1));
  reg_module u_reg_t0_15_d5 (.clk(clk), .input_share0(d4_t0_15_s0), .input_share1(d4_t0_15_s1), .output_share0(d5_t0_15_s0), .output_share1(d5_t0_15_s1));
  reg_module u_reg_t0_16_d5 (.clk(clk), .input_share0(d4_t0_16_s0), .input_share1(d4_t0_16_s1), .output_share0(d5_t0_16_s0), .output_share1(d5_t0_16_s1));
  reg_module u_reg_t0_17_d5 (.clk(clk), .input_share0(d4_t0_17_s0), .input_share1(d4_t0_17_s1), .output_share0(d5_t0_17_s0), .output_share1(d5_t0_17_s1));
  reg_module u_reg_t0_18_d5 (.clk(clk), .input_share0(d4_t0_18_s0), .input_share1(d4_t0_18_s1), .output_share0(d5_t0_18_s0), .output_share1(d5_t0_18_s1));
  reg_module u_reg_t0_19_d5 (.clk(clk), .input_share0(d4_t0_19_s0), .input_share1(d4_t0_19_s1), .output_share0(d5_t0_19_s0), .output_share1(d5_t0_19_s1));
  reg_module u_reg_t0_20_d5 (.clk(clk), .input_share0(d4_t0_20_s0), .input_share1(d4_t0_20_s1), .output_share0(d5_t0_20_s0), .output_share1(d5_t0_20_s1));
  reg_module u_reg_t0_21_d5 (.clk(clk), .input_share0(d4_t0_21_s0), .input_share1(d4_t0_21_s1), .output_share0(d5_t0_21_s0), .output_share1(d5_t0_21_s1));
  reg_module u_reg_t0_22_d5 (.clk(clk), .input_share0(d4_t0_22_s0), .input_share1(d4_t0_22_s1), .output_share0(d5_t0_22_s0), .output_share1(d5_t0_22_s1));
  reg_module u_reg_t0_23_d5 (.clk(clk), .input_share0(d4_t0_23_s0), .input_share1(d4_t0_23_s1), .output_share0(d5_t0_23_s0), .output_share1(d5_t0_23_s1));
  reg_module u_reg_t0_24_d5 (.clk(clk), .input_share0(d4_t0_24_s0), .input_share1(d4_t0_24_s1), .output_share0(d5_t0_24_s0), .output_share1(d5_t0_24_s1));
  reg_module u_reg_t0_25_d5 (.clk(clk), .input_share0(d4_t0_25_s0), .input_share1(d4_t0_25_s1), .output_share0(d5_t0_25_s0), .output_share1(d5_t0_25_s1));
  reg_module u_reg_t0_26_d5 (.clk(clk), .input_share0(d4_t0_26_s0), .input_share1(d4_t0_26_s1), .output_share0(d5_t0_26_s0), .output_share1(d5_t0_26_s1));
  reg_module u_reg_t0_27_d5 (.clk(clk), .input_share0(d4_t0_27_s0), .input_share1(d4_t0_27_s1), .output_share0(d5_t0_27_s0), .output_share1(d5_t0_27_s1));
  reg_module u_reg_t0_28_d5 (.clk(clk), .input_share0(d4_t0_28_s0), .input_share1(d4_t0_28_s1), .output_share0(d5_t0_28_s0), .output_share1(d5_t0_28_s1));
  reg_module u_reg_t0_29_d5 (.clk(clk), .input_share0(d4_t0_29_s0), .input_share1(d4_t0_29_s1), .output_share0(d5_t0_29_s0), .output_share1(d5_t0_29_s1));
  reg_module u_reg_t0_30_d5 (.clk(clk), .input_share0(d4_t0_30_s0), .input_share1(d4_t0_30_s1), .output_share0(d5_t0_30_s0), .output_share1(d5_t0_30_s1));
  reg_module u_reg_t0_31_d5 (.clk(clk), .input_share0(d4_t0_31_s0), .input_share1(d4_t0_31_s1), .output_share0(d5_t0_31_s0), .output_share1(d5_t0_31_s1));
  reg_module u_reg_t0_5_d5 (.clk(clk), .input_share0(d4_t0_5_s0), .input_share1(d4_t0_5_s1), .output_share0(d5_t0_5_s0), .output_share1(d5_t0_5_s1));
  reg_module u_reg_t0_6_d5 (.clk(clk), .input_share0(d4_t0_6_s0), .input_share1(d4_t0_6_s1), .output_share0(d5_t0_6_s0), .output_share1(d5_t0_6_s1));
  reg_module u_reg_t0_7_d5 (.clk(clk), .input_share0(d4_t0_7_s0), .input_share1(d4_t0_7_s1), .output_share0(d5_t0_7_s0), .output_share1(d5_t0_7_s1));
  reg_module u_reg_t0_8_d5 (.clk(clk), .input_share0(d4_t0_8_s0), .input_share1(d4_t0_8_s1), .output_share0(d5_t0_8_s0), .output_share1(d5_t0_8_s1));
  reg_module u_reg_t0_9_d5 (.clk(clk), .input_share0(d4_t0_9_s0), .input_share1(d4_t0_9_s1), .output_share0(d5_t0_9_s0), .output_share1(d5_t0_9_s1));
  xor_module u_xor_c5_d5 (.x_share0(d5_i4_s0), .x_share1(d5_i4_s1), .y_share0(d5_t2_4_s0), .y_share1(d5_t2_4_s1), .z_share0(d5_c5_s0), .z_share1(d5_c5_s1));
  xor_module u_xor_o5_d5 (.x_share0(d5_t0_5_s0), .x_share1(d5_t0_5_s1), .y_share0(d5_c5_s0), .y_share1(d5_c5_s1), .z_share0(d5_o5_s0), .z_share1(d5_o5_s1));
  xor_module u_xor_t1_5_d5 (.x_share0(d5_i5_s0), .x_share1(d5_i5_s1), .y_share0(d5_c5_s0), .y_share1(d5_c5_s1), .z_share0(d5_t1_5_s0), .z_share1(d5_t1_5_s1));
  and_module u_and_t2_4_d5 (.clk(clk), .x_share0(d4_t0_4_s0), .x_share1(d4_t0_4_s1), .y_share0(d4_t1_4_s0), .y_share1(d4_t1_4_s1), .rand(r_t2_4), .z_share0(d5_t2_4_s0), .z_share1(d5_t2_4_s1));
  assign r_t2_4 = stage5_share0[2];
  reg_module u_reg_i10_d6 (.clk(clk), .input_share0(d5_i10_s0), .input_share1(d5_i10_s1), .output_share0(d6_i10_s0), .output_share1(d6_i10_s1));
  reg_module u_reg_i11_d6 (.clk(clk), .input_share0(d5_i11_s0), .input_share1(d5_i11_s1), .output_share0(d6_i11_s0), .output_share1(d6_i11_s1));
  reg_module u_reg_i12_d6 (.clk(clk), .input_share0(d5_i12_s0), .input_share1(d5_i12_s1), .output_share0(d6_i12_s0), .output_share1(d6_i12_s1));
  reg_module u_reg_i13_d6 (.clk(clk), .input_share0(d5_i13_s0), .input_share1(d5_i13_s1), .output_share0(d6_i13_s0), .output_share1(d6_i13_s1));
  reg_module u_reg_i14_d6 (.clk(clk), .input_share0(d5_i14_s0), .input_share1(d5_i14_s1), .output_share0(d6_i14_s0), .output_share1(d6_i14_s1));
  reg_module u_reg_i15_d6 (.clk(clk), .input_share0(d5_i15_s0), .input_share1(d5_i15_s1), .output_share0(d6_i15_s0), .output_share1(d6_i15_s1));
  reg_module u_reg_i16_d6 (.clk(clk), .input_share0(d5_i16_s0), .input_share1(d5_i16_s1), .output_share0(d6_i16_s0), .output_share1(d6_i16_s1));
  reg_module u_reg_i17_d6 (.clk(clk), .input_share0(d5_i17_s0), .input_share1(d5_i17_s1), .output_share0(d6_i17_s0), .output_share1(d6_i17_s1));
  reg_module u_reg_i18_d6 (.clk(clk), .input_share0(d5_i18_s0), .input_share1(d5_i18_s1), .output_share0(d6_i18_s0), .output_share1(d6_i18_s1));
  reg_module u_reg_i19_d6 (.clk(clk), .input_share0(d5_i19_s0), .input_share1(d5_i19_s1), .output_share0(d6_i19_s0), .output_share1(d6_i19_s1));
  reg_module u_reg_i20_d6 (.clk(clk), .input_share0(d5_i20_s0), .input_share1(d5_i20_s1), .output_share0(d6_i20_s0), .output_share1(d6_i20_s1));
  reg_module u_reg_i21_d6 (.clk(clk), .input_share0(d5_i21_s0), .input_share1(d5_i21_s1), .output_share0(d6_i21_s0), .output_share1(d6_i21_s1));
  reg_module u_reg_i22_d6 (.clk(clk), .input_share0(d5_i22_s0), .input_share1(d5_i22_s1), .output_share0(d6_i22_s0), .output_share1(d6_i22_s1));
  reg_module u_reg_i23_d6 (.clk(clk), .input_share0(d5_i23_s0), .input_share1(d5_i23_s1), .output_share0(d6_i23_s0), .output_share1(d6_i23_s1));
  reg_module u_reg_i24_d6 (.clk(clk), .input_share0(d5_i24_s0), .input_share1(d5_i24_s1), .output_share0(d6_i24_s0), .output_share1(d6_i24_s1));
  reg_module u_reg_i25_d6 (.clk(clk), .input_share0(d5_i25_s0), .input_share1(d5_i25_s1), .output_share0(d6_i25_s0), .output_share1(d6_i25_s1));
  reg_module u_reg_i26_d6 (.clk(clk), .input_share0(d5_i26_s0), .input_share1(d5_i26_s1), .output_share0(d6_i26_s0), .output_share1(d6_i26_s1));
  reg_module u_reg_i27_d6 (.clk(clk), .input_share0(d5_i27_s0), .input_share1(d5_i27_s1), .output_share0(d6_i27_s0), .output_share1(d6_i27_s1));
  reg_module u_reg_i28_d6 (.clk(clk), .input_share0(d5_i28_s0), .input_share1(d5_i28_s1), .output_share0(d6_i28_s0), .output_share1(d6_i28_s1));
  reg_module u_reg_i29_d6 (.clk(clk), .input_share0(d5_i29_s0), .input_share1(d5_i29_s1), .output_share0(d6_i29_s0), .output_share1(d6_i29_s1));
  reg_module u_reg_i30_d6 (.clk(clk), .input_share0(d5_i30_s0), .input_share1(d5_i30_s1), .output_share0(d6_i30_s0), .output_share1(d6_i30_s1));
  reg_module u_reg_i5_d6 (.clk(clk), .input_share0(d5_i5_s0), .input_share1(d5_i5_s1), .output_share0(d6_i5_s0), .output_share1(d6_i5_s1));
  reg_module u_reg_i6_d6 (.clk(clk), .input_share0(d5_i6_s0), .input_share1(d5_i6_s1), .output_share0(d6_i6_s0), .output_share1(d6_i6_s1));
  reg_module u_reg_i7_d6 (.clk(clk), .input_share0(d5_i7_s0), .input_share1(d5_i7_s1), .output_share0(d6_i7_s0), .output_share1(d6_i7_s1));
  reg_module u_reg_i8_d6 (.clk(clk), .input_share0(d5_i8_s0), .input_share1(d5_i8_s1), .output_share0(d6_i8_s0), .output_share1(d6_i8_s1));
  reg_module u_reg_i9_d6 (.clk(clk), .input_share0(d5_i9_s0), .input_share1(d5_i9_s1), .output_share0(d6_i9_s0), .output_share1(d6_i9_s1));
  reg_module u_reg_t0_10_d6 (.clk(clk), .input_share0(d5_t0_10_s0), .input_share1(d5_t0_10_s1), .output_share0(d6_t0_10_s0), .output_share1(d6_t0_10_s1));
  reg_module u_reg_t0_11_d6 (.clk(clk), .input_share0(d5_t0_11_s0), .input_share1(d5_t0_11_s1), .output_share0(d6_t0_11_s0), .output_share1(d6_t0_11_s1));
  reg_module u_reg_t0_12_d6 (.clk(clk), .input_share0(d5_t0_12_s0), .input_share1(d5_t0_12_s1), .output_share0(d6_t0_12_s0), .output_share1(d6_t0_12_s1));
  reg_module u_reg_t0_13_d6 (.clk(clk), .input_share0(d5_t0_13_s0), .input_share1(d5_t0_13_s1), .output_share0(d6_t0_13_s0), .output_share1(d6_t0_13_s1));
  reg_module u_reg_t0_14_d6 (.clk(clk), .input_share0(d5_t0_14_s0), .input_share1(d5_t0_14_s1), .output_share0(d6_t0_14_s0), .output_share1(d6_t0_14_s1));
  reg_module u_reg_t0_15_d6 (.clk(clk), .input_share0(d5_t0_15_s0), .input_share1(d5_t0_15_s1), .output_share0(d6_t0_15_s0), .output_share1(d6_t0_15_s1));
  reg_module u_reg_t0_16_d6 (.clk(clk), .input_share0(d5_t0_16_s0), .input_share1(d5_t0_16_s1), .output_share0(d6_t0_16_s0), .output_share1(d6_t0_16_s1));
  reg_module u_reg_t0_17_d6 (.clk(clk), .input_share0(d5_t0_17_s0), .input_share1(d5_t0_17_s1), .output_share0(d6_t0_17_s0), .output_share1(d6_t0_17_s1));
  reg_module u_reg_t0_18_d6 (.clk(clk), .input_share0(d5_t0_18_s0), .input_share1(d5_t0_18_s1), .output_share0(d6_t0_18_s0), .output_share1(d6_t0_18_s1));
  reg_module u_reg_t0_19_d6 (.clk(clk), .input_share0(d5_t0_19_s0), .input_share1(d5_t0_19_s1), .output_share0(d6_t0_19_s0), .output_share1(d6_t0_19_s1));
  reg_module u_reg_t0_20_d6 (.clk(clk), .input_share0(d5_t0_20_s0), .input_share1(d5_t0_20_s1), .output_share0(d6_t0_20_s0), .output_share1(d6_t0_20_s1));
  reg_module u_reg_t0_21_d6 (.clk(clk), .input_share0(d5_t0_21_s0), .input_share1(d5_t0_21_s1), .output_share0(d6_t0_21_s0), .output_share1(d6_t0_21_s1));
  reg_module u_reg_t0_22_d6 (.clk(clk), .input_share0(d5_t0_22_s0), .input_share1(d5_t0_22_s1), .output_share0(d6_t0_22_s0), .output_share1(d6_t0_22_s1));
  reg_module u_reg_t0_23_d6 (.clk(clk), .input_share0(d5_t0_23_s0), .input_share1(d5_t0_23_s1), .output_share0(d6_t0_23_s0), .output_share1(d6_t0_23_s1));
  reg_module u_reg_t0_24_d6 (.clk(clk), .input_share0(d5_t0_24_s0), .input_share1(d5_t0_24_s1), .output_share0(d6_t0_24_s0), .output_share1(d6_t0_24_s1));
  reg_module u_reg_t0_25_d6 (.clk(clk), .input_share0(d5_t0_25_s0), .input_share1(d5_t0_25_s1), .output_share0(d6_t0_25_s0), .output_share1(d6_t0_25_s1));
  reg_module u_reg_t0_26_d6 (.clk(clk), .input_share0(d5_t0_26_s0), .input_share1(d5_t0_26_s1), .output_share0(d6_t0_26_s0), .output_share1(d6_t0_26_s1));
  reg_module u_reg_t0_27_d6 (.clk(clk), .input_share0(d5_t0_27_s0), .input_share1(d5_t0_27_s1), .output_share0(d6_t0_27_s0), .output_share1(d6_t0_27_s1));
  reg_module u_reg_t0_28_d6 (.clk(clk), .input_share0(d5_t0_28_s0), .input_share1(d5_t0_28_s1), .output_share0(d6_t0_28_s0), .output_share1(d6_t0_28_s1));
  reg_module u_reg_t0_29_d6 (.clk(clk), .input_share0(d5_t0_29_s0), .input_share1(d5_t0_29_s1), .output_share0(d6_t0_29_s0), .output_share1(d6_t0_29_s1));
  reg_module u_reg_t0_30_d6 (.clk(clk), .input_share0(d5_t0_30_s0), .input_share1(d5_t0_30_s1), .output_share0(d6_t0_30_s0), .output_share1(d6_t0_30_s1));
  reg_module u_reg_t0_31_d6 (.clk(clk), .input_share0(d5_t0_31_s0), .input_share1(d5_t0_31_s1), .output_share0(d6_t0_31_s0), .output_share1(d6_t0_31_s1));
  reg_module u_reg_t0_6_d6 (.clk(clk), .input_share0(d5_t0_6_s0), .input_share1(d5_t0_6_s1), .output_share0(d6_t0_6_s0), .output_share1(d6_t0_6_s1));
  reg_module u_reg_t0_7_d6 (.clk(clk), .input_share0(d5_t0_7_s0), .input_share1(d5_t0_7_s1), .output_share0(d6_t0_7_s0), .output_share1(d6_t0_7_s1));
  reg_module u_reg_t0_8_d6 (.clk(clk), .input_share0(d5_t0_8_s0), .input_share1(d5_t0_8_s1), .output_share0(d6_t0_8_s0), .output_share1(d6_t0_8_s1));
  reg_module u_reg_t0_9_d6 (.clk(clk), .input_share0(d5_t0_9_s0), .input_share1(d5_t0_9_s1), .output_share0(d6_t0_9_s0), .output_share1(d6_t0_9_s1));
  xor_module u_xor_c6_d6 (.x_share0(d6_i5_s0), .x_share1(d6_i5_s1), .y_share0(d6_t2_5_s0), .y_share1(d6_t2_5_s1), .z_share0(d6_c6_s0), .z_share1(d6_c6_s1));
  xor_module u_xor_o6_d6 (.x_share0(d6_t0_6_s0), .x_share1(d6_t0_6_s1), .y_share0(d6_c6_s0), .y_share1(d6_c6_s1), .z_share0(d6_o6_s0), .z_share1(d6_o6_s1));
  xor_module u_xor_t1_6_d6 (.x_share0(d6_i6_s0), .x_share1(d6_i6_s1), .y_share0(d6_c6_s0), .y_share1(d6_c6_s1), .z_share0(d6_t1_6_s0), .z_share1(d6_t1_6_s1));
  and_module u_and_t2_5_d6 (.clk(clk), .x_share0(d5_t0_5_s0), .x_share1(d5_t0_5_s1), .y_share0(d5_t1_5_s0), .y_share1(d5_t1_5_s1), .rand(r_t2_5), .z_share0(d6_t2_5_s0), .z_share1(d6_t2_5_s1));
  assign r_t2_5 = stage6_share0[0];
  reg_module u_reg_i10_d7 (.clk(clk), .input_share0(d6_i10_s0), .input_share1(d6_i10_s1), .output_share0(d7_i10_s0), .output_share1(d7_i10_s1));
  reg_module u_reg_i11_d7 (.clk(clk), .input_share0(d6_i11_s0), .input_share1(d6_i11_s1), .output_share0(d7_i11_s0), .output_share1(d7_i11_s1));
  reg_module u_reg_i12_d7 (.clk(clk), .input_share0(d6_i12_s0), .input_share1(d6_i12_s1), .output_share0(d7_i12_s0), .output_share1(d7_i12_s1));
  reg_module u_reg_i13_d7 (.clk(clk), .input_share0(d6_i13_s0), .input_share1(d6_i13_s1), .output_share0(d7_i13_s0), .output_share1(d7_i13_s1));
  reg_module u_reg_i14_d7 (.clk(clk), .input_share0(d6_i14_s0), .input_share1(d6_i14_s1), .output_share0(d7_i14_s0), .output_share1(d7_i14_s1));
  reg_module u_reg_i15_d7 (.clk(clk), .input_share0(d6_i15_s0), .input_share1(d6_i15_s1), .output_share0(d7_i15_s0), .output_share1(d7_i15_s1));
  reg_module u_reg_i16_d7 (.clk(clk), .input_share0(d6_i16_s0), .input_share1(d6_i16_s1), .output_share0(d7_i16_s0), .output_share1(d7_i16_s1));
  reg_module u_reg_i17_d7 (.clk(clk), .input_share0(d6_i17_s0), .input_share1(d6_i17_s1), .output_share0(d7_i17_s0), .output_share1(d7_i17_s1));
  reg_module u_reg_i18_d7 (.clk(clk), .input_share0(d6_i18_s0), .input_share1(d6_i18_s1), .output_share0(d7_i18_s0), .output_share1(d7_i18_s1));
  reg_module u_reg_i19_d7 (.clk(clk), .input_share0(d6_i19_s0), .input_share1(d6_i19_s1), .output_share0(d7_i19_s0), .output_share1(d7_i19_s1));
  reg_module u_reg_i20_d7 (.clk(clk), .input_share0(d6_i20_s0), .input_share1(d6_i20_s1), .output_share0(d7_i20_s0), .output_share1(d7_i20_s1));
  reg_module u_reg_i21_d7 (.clk(clk), .input_share0(d6_i21_s0), .input_share1(d6_i21_s1), .output_share0(d7_i21_s0), .output_share1(d7_i21_s1));
  reg_module u_reg_i22_d7 (.clk(clk), .input_share0(d6_i22_s0), .input_share1(d6_i22_s1), .output_share0(d7_i22_s0), .output_share1(d7_i22_s1));
  reg_module u_reg_i23_d7 (.clk(clk), .input_share0(d6_i23_s0), .input_share1(d6_i23_s1), .output_share0(d7_i23_s0), .output_share1(d7_i23_s1));
  reg_module u_reg_i24_d7 (.clk(clk), .input_share0(d6_i24_s0), .input_share1(d6_i24_s1), .output_share0(d7_i24_s0), .output_share1(d7_i24_s1));
  reg_module u_reg_i25_d7 (.clk(clk), .input_share0(d6_i25_s0), .input_share1(d6_i25_s1), .output_share0(d7_i25_s0), .output_share1(d7_i25_s1));
  reg_module u_reg_i26_d7 (.clk(clk), .input_share0(d6_i26_s0), .input_share1(d6_i26_s1), .output_share0(d7_i26_s0), .output_share1(d7_i26_s1));
  reg_module u_reg_i27_d7 (.clk(clk), .input_share0(d6_i27_s0), .input_share1(d6_i27_s1), .output_share0(d7_i27_s0), .output_share1(d7_i27_s1));
  reg_module u_reg_i28_d7 (.clk(clk), .input_share0(d6_i28_s0), .input_share1(d6_i28_s1), .output_share0(d7_i28_s0), .output_share1(d7_i28_s1));
  reg_module u_reg_i29_d7 (.clk(clk), .input_share0(d6_i29_s0), .input_share1(d6_i29_s1), .output_share0(d7_i29_s0), .output_share1(d7_i29_s1));
  reg_module u_reg_i30_d7 (.clk(clk), .input_share0(d6_i30_s0), .input_share1(d6_i30_s1), .output_share0(d7_i30_s0), .output_share1(d7_i30_s1));
  reg_module u_reg_i6_d7 (.clk(clk), .input_share0(d6_i6_s0), .input_share1(d6_i6_s1), .output_share0(d7_i6_s0), .output_share1(d7_i6_s1));
  reg_module u_reg_i7_d7 (.clk(clk), .input_share0(d6_i7_s0), .input_share1(d6_i7_s1), .output_share0(d7_i7_s0), .output_share1(d7_i7_s1));
  reg_module u_reg_i8_d7 (.clk(clk), .input_share0(d6_i8_s0), .input_share1(d6_i8_s1), .output_share0(d7_i8_s0), .output_share1(d7_i8_s1));
  reg_module u_reg_i9_d7 (.clk(clk), .input_share0(d6_i9_s0), .input_share1(d6_i9_s1), .output_share0(d7_i9_s0), .output_share1(d7_i9_s1));
  reg_module u_reg_t0_10_d7 (.clk(clk), .input_share0(d6_t0_10_s0), .input_share1(d6_t0_10_s1), .output_share0(d7_t0_10_s0), .output_share1(d7_t0_10_s1));
  reg_module u_reg_t0_11_d7 (.clk(clk), .input_share0(d6_t0_11_s0), .input_share1(d6_t0_11_s1), .output_share0(d7_t0_11_s0), .output_share1(d7_t0_11_s1));
  reg_module u_reg_t0_12_d7 (.clk(clk), .input_share0(d6_t0_12_s0), .input_share1(d6_t0_12_s1), .output_share0(d7_t0_12_s0), .output_share1(d7_t0_12_s1));
  reg_module u_reg_t0_13_d7 (.clk(clk), .input_share0(d6_t0_13_s0), .input_share1(d6_t0_13_s1), .output_share0(d7_t0_13_s0), .output_share1(d7_t0_13_s1));
  reg_module u_reg_t0_14_d7 (.clk(clk), .input_share0(d6_t0_14_s0), .input_share1(d6_t0_14_s1), .output_share0(d7_t0_14_s0), .output_share1(d7_t0_14_s1));
  reg_module u_reg_t0_15_d7 (.clk(clk), .input_share0(d6_t0_15_s0), .input_share1(d6_t0_15_s1), .output_share0(d7_t0_15_s0), .output_share1(d7_t0_15_s1));
  reg_module u_reg_t0_16_d7 (.clk(clk), .input_share0(d6_t0_16_s0), .input_share1(d6_t0_16_s1), .output_share0(d7_t0_16_s0), .output_share1(d7_t0_16_s1));
  reg_module u_reg_t0_17_d7 (.clk(clk), .input_share0(d6_t0_17_s0), .input_share1(d6_t0_17_s1), .output_share0(d7_t0_17_s0), .output_share1(d7_t0_17_s1));
  reg_module u_reg_t0_18_d7 (.clk(clk), .input_share0(d6_t0_18_s0), .input_share1(d6_t0_18_s1), .output_share0(d7_t0_18_s0), .output_share1(d7_t0_18_s1));
  reg_module u_reg_t0_19_d7 (.clk(clk), .input_share0(d6_t0_19_s0), .input_share1(d6_t0_19_s1), .output_share0(d7_t0_19_s0), .output_share1(d7_t0_19_s1));
  reg_module u_reg_t0_20_d7 (.clk(clk), .input_share0(d6_t0_20_s0), .input_share1(d6_t0_20_s1), .output_share0(d7_t0_20_s0), .output_share1(d7_t0_20_s1));
  reg_module u_reg_t0_21_d7 (.clk(clk), .input_share0(d6_t0_21_s0), .input_share1(d6_t0_21_s1), .output_share0(d7_t0_21_s0), .output_share1(d7_t0_21_s1));
  reg_module u_reg_t0_22_d7 (.clk(clk), .input_share0(d6_t0_22_s0), .input_share1(d6_t0_22_s1), .output_share0(d7_t0_22_s0), .output_share1(d7_t0_22_s1));
  reg_module u_reg_t0_23_d7 (.clk(clk), .input_share0(d6_t0_23_s0), .input_share1(d6_t0_23_s1), .output_share0(d7_t0_23_s0), .output_share1(d7_t0_23_s1));
  reg_module u_reg_t0_24_d7 (.clk(clk), .input_share0(d6_t0_24_s0), .input_share1(d6_t0_24_s1), .output_share0(d7_t0_24_s0), .output_share1(d7_t0_24_s1));
  reg_module u_reg_t0_25_d7 (.clk(clk), .input_share0(d6_t0_25_s0), .input_share1(d6_t0_25_s1), .output_share0(d7_t0_25_s0), .output_share1(d7_t0_25_s1));
  reg_module u_reg_t0_26_d7 (.clk(clk), .input_share0(d6_t0_26_s0), .input_share1(d6_t0_26_s1), .output_share0(d7_t0_26_s0), .output_share1(d7_t0_26_s1));
  reg_module u_reg_t0_27_d7 (.clk(clk), .input_share0(d6_t0_27_s0), .input_share1(d6_t0_27_s1), .output_share0(d7_t0_27_s0), .output_share1(d7_t0_27_s1));
  reg_module u_reg_t0_28_d7 (.clk(clk), .input_share0(d6_t0_28_s0), .input_share1(d6_t0_28_s1), .output_share0(d7_t0_28_s0), .output_share1(d7_t0_28_s1));
  reg_module u_reg_t0_29_d7 (.clk(clk), .input_share0(d6_t0_29_s0), .input_share1(d6_t0_29_s1), .output_share0(d7_t0_29_s0), .output_share1(d7_t0_29_s1));
  reg_module u_reg_t0_30_d7 (.clk(clk), .input_share0(d6_t0_30_s0), .input_share1(d6_t0_30_s1), .output_share0(d7_t0_30_s0), .output_share1(d7_t0_30_s1));
  reg_module u_reg_t0_31_d7 (.clk(clk), .input_share0(d6_t0_31_s0), .input_share1(d6_t0_31_s1), .output_share0(d7_t0_31_s0), .output_share1(d7_t0_31_s1));
  reg_module u_reg_t0_7_d7 (.clk(clk), .input_share0(d6_t0_7_s0), .input_share1(d6_t0_7_s1), .output_share0(d7_t0_7_s0), .output_share1(d7_t0_7_s1));
  reg_module u_reg_t0_8_d7 (.clk(clk), .input_share0(d6_t0_8_s0), .input_share1(d6_t0_8_s1), .output_share0(d7_t0_8_s0), .output_share1(d7_t0_8_s1));
  reg_module u_reg_t0_9_d7 (.clk(clk), .input_share0(d6_t0_9_s0), .input_share1(d6_t0_9_s1), .output_share0(d7_t0_9_s0), .output_share1(d7_t0_9_s1));
  xor_module u_xor_c7_d7 (.x_share0(d7_i6_s0), .x_share1(d7_i6_s1), .y_share0(d7_t2_6_s0), .y_share1(d7_t2_6_s1), .z_share0(d7_c7_s0), .z_share1(d7_c7_s1));
  xor_module u_xor_o7_d7 (.x_share0(d7_t0_7_s0), .x_share1(d7_t0_7_s1), .y_share0(d7_c7_s0), .y_share1(d7_c7_s1), .z_share0(d7_o7_s0), .z_share1(d7_o7_s1));
  xor_module u_xor_t1_7_d7 (.x_share0(d7_i7_s0), .x_share1(d7_i7_s1), .y_share0(d7_c7_s0), .y_share1(d7_c7_s1), .z_share0(d7_t1_7_s0), .z_share1(d7_t1_7_s1));
  and_module u_and_t2_6_d7 (.clk(clk), .x_share0(d6_t0_6_s0), .x_share1(d6_t0_6_s1), .y_share0(d6_t1_6_s0), .y_share1(d6_t1_6_s1), .rand(r_t2_6), .z_share0(d7_t2_6_s0), .z_share1(d7_t2_6_s1));
  assign r_t2_6 = stage7_share0[1];
  reg_module u_reg_i10_d8 (.clk(clk), .input_share0(d7_i10_s0), .input_share1(d7_i10_s1), .output_share0(d8_i10_s0), .output_share1(d8_i10_s1));
  reg_module u_reg_i11_d8 (.clk(clk), .input_share0(d7_i11_s0), .input_share1(d7_i11_s1), .output_share0(d8_i11_s0), .output_share1(d8_i11_s1));
  reg_module u_reg_i12_d8 (.clk(clk), .input_share0(d7_i12_s0), .input_share1(d7_i12_s1), .output_share0(d8_i12_s0), .output_share1(d8_i12_s1));
  reg_module u_reg_i13_d8 (.clk(clk), .input_share0(d7_i13_s0), .input_share1(d7_i13_s1), .output_share0(d8_i13_s0), .output_share1(d8_i13_s1));
  reg_module u_reg_i14_d8 (.clk(clk), .input_share0(d7_i14_s0), .input_share1(d7_i14_s1), .output_share0(d8_i14_s0), .output_share1(d8_i14_s1));
  reg_module u_reg_i15_d8 (.clk(clk), .input_share0(d7_i15_s0), .input_share1(d7_i15_s1), .output_share0(d8_i15_s0), .output_share1(d8_i15_s1));
  reg_module u_reg_i16_d8 (.clk(clk), .input_share0(d7_i16_s0), .input_share1(d7_i16_s1), .output_share0(d8_i16_s0), .output_share1(d8_i16_s1));
  reg_module u_reg_i17_d8 (.clk(clk), .input_share0(d7_i17_s0), .input_share1(d7_i17_s1), .output_share0(d8_i17_s0), .output_share1(d8_i17_s1));
  reg_module u_reg_i18_d8 (.clk(clk), .input_share0(d7_i18_s0), .input_share1(d7_i18_s1), .output_share0(d8_i18_s0), .output_share1(d8_i18_s1));
  reg_module u_reg_i19_d8 (.clk(clk), .input_share0(d7_i19_s0), .input_share1(d7_i19_s1), .output_share0(d8_i19_s0), .output_share1(d8_i19_s1));
  reg_module u_reg_i20_d8 (.clk(clk), .input_share0(d7_i20_s0), .input_share1(d7_i20_s1), .output_share0(d8_i20_s0), .output_share1(d8_i20_s1));
  reg_module u_reg_i21_d8 (.clk(clk), .input_share0(d7_i21_s0), .input_share1(d7_i21_s1), .output_share0(d8_i21_s0), .output_share1(d8_i21_s1));
  reg_module u_reg_i22_d8 (.clk(clk), .input_share0(d7_i22_s0), .input_share1(d7_i22_s1), .output_share0(d8_i22_s0), .output_share1(d8_i22_s1));
  reg_module u_reg_i23_d8 (.clk(clk), .input_share0(d7_i23_s0), .input_share1(d7_i23_s1), .output_share0(d8_i23_s0), .output_share1(d8_i23_s1));
  reg_module u_reg_i24_d8 (.clk(clk), .input_share0(d7_i24_s0), .input_share1(d7_i24_s1), .output_share0(d8_i24_s0), .output_share1(d8_i24_s1));
  reg_module u_reg_i25_d8 (.clk(clk), .input_share0(d7_i25_s0), .input_share1(d7_i25_s1), .output_share0(d8_i25_s0), .output_share1(d8_i25_s1));
  reg_module u_reg_i26_d8 (.clk(clk), .input_share0(d7_i26_s0), .input_share1(d7_i26_s1), .output_share0(d8_i26_s0), .output_share1(d8_i26_s1));
  reg_module u_reg_i27_d8 (.clk(clk), .input_share0(d7_i27_s0), .input_share1(d7_i27_s1), .output_share0(d8_i27_s0), .output_share1(d8_i27_s1));
  reg_module u_reg_i28_d8 (.clk(clk), .input_share0(d7_i28_s0), .input_share1(d7_i28_s1), .output_share0(d8_i28_s0), .output_share1(d8_i28_s1));
  reg_module u_reg_i29_d8 (.clk(clk), .input_share0(d7_i29_s0), .input_share1(d7_i29_s1), .output_share0(d8_i29_s0), .output_share1(d8_i29_s1));
  reg_module u_reg_i30_d8 (.clk(clk), .input_share0(d7_i30_s0), .input_share1(d7_i30_s1), .output_share0(d8_i30_s0), .output_share1(d8_i30_s1));
  reg_module u_reg_i7_d8 (.clk(clk), .input_share0(d7_i7_s0), .input_share1(d7_i7_s1), .output_share0(d8_i7_s0), .output_share1(d8_i7_s1));
  reg_module u_reg_i8_d8 (.clk(clk), .input_share0(d7_i8_s0), .input_share1(d7_i8_s1), .output_share0(d8_i8_s0), .output_share1(d8_i8_s1));
  reg_module u_reg_i9_d8 (.clk(clk), .input_share0(d7_i9_s0), .input_share1(d7_i9_s1), .output_share0(d8_i9_s0), .output_share1(d8_i9_s1));
  reg_module u_reg_t0_10_d8 (.clk(clk), .input_share0(d7_t0_10_s0), .input_share1(d7_t0_10_s1), .output_share0(d8_t0_10_s0), .output_share1(d8_t0_10_s1));
  reg_module u_reg_t0_11_d8 (.clk(clk), .input_share0(d7_t0_11_s0), .input_share1(d7_t0_11_s1), .output_share0(d8_t0_11_s0), .output_share1(d8_t0_11_s1));
  reg_module u_reg_t0_12_d8 (.clk(clk), .input_share0(d7_t0_12_s0), .input_share1(d7_t0_12_s1), .output_share0(d8_t0_12_s0), .output_share1(d8_t0_12_s1));
  reg_module u_reg_t0_13_d8 (.clk(clk), .input_share0(d7_t0_13_s0), .input_share1(d7_t0_13_s1), .output_share0(d8_t0_13_s0), .output_share1(d8_t0_13_s1));
  reg_module u_reg_t0_14_d8 (.clk(clk), .input_share0(d7_t0_14_s0), .input_share1(d7_t0_14_s1), .output_share0(d8_t0_14_s0), .output_share1(d8_t0_14_s1));
  reg_module u_reg_t0_15_d8 (.clk(clk), .input_share0(d7_t0_15_s0), .input_share1(d7_t0_15_s1), .output_share0(d8_t0_15_s0), .output_share1(d8_t0_15_s1));
  reg_module u_reg_t0_16_d8 (.clk(clk), .input_share0(d7_t0_16_s0), .input_share1(d7_t0_16_s1), .output_share0(d8_t0_16_s0), .output_share1(d8_t0_16_s1));
  reg_module u_reg_t0_17_d8 (.clk(clk), .input_share0(d7_t0_17_s0), .input_share1(d7_t0_17_s1), .output_share0(d8_t0_17_s0), .output_share1(d8_t0_17_s1));
  reg_module u_reg_t0_18_d8 (.clk(clk), .input_share0(d7_t0_18_s0), .input_share1(d7_t0_18_s1), .output_share0(d8_t0_18_s0), .output_share1(d8_t0_18_s1));
  reg_module u_reg_t0_19_d8 (.clk(clk), .input_share0(d7_t0_19_s0), .input_share1(d7_t0_19_s1), .output_share0(d8_t0_19_s0), .output_share1(d8_t0_19_s1));
  reg_module u_reg_t0_20_d8 (.clk(clk), .input_share0(d7_t0_20_s0), .input_share1(d7_t0_20_s1), .output_share0(d8_t0_20_s0), .output_share1(d8_t0_20_s1));
  reg_module u_reg_t0_21_d8 (.clk(clk), .input_share0(d7_t0_21_s0), .input_share1(d7_t0_21_s1), .output_share0(d8_t0_21_s0), .output_share1(d8_t0_21_s1));
  reg_module u_reg_t0_22_d8 (.clk(clk), .input_share0(d7_t0_22_s0), .input_share1(d7_t0_22_s1), .output_share0(d8_t0_22_s0), .output_share1(d8_t0_22_s1));
  reg_module u_reg_t0_23_d8 (.clk(clk), .input_share0(d7_t0_23_s0), .input_share1(d7_t0_23_s1), .output_share0(d8_t0_23_s0), .output_share1(d8_t0_23_s1));
  reg_module u_reg_t0_24_d8 (.clk(clk), .input_share0(d7_t0_24_s0), .input_share1(d7_t0_24_s1), .output_share0(d8_t0_24_s0), .output_share1(d8_t0_24_s1));
  reg_module u_reg_t0_25_d8 (.clk(clk), .input_share0(d7_t0_25_s0), .input_share1(d7_t0_25_s1), .output_share0(d8_t0_25_s0), .output_share1(d8_t0_25_s1));
  reg_module u_reg_t0_26_d8 (.clk(clk), .input_share0(d7_t0_26_s0), .input_share1(d7_t0_26_s1), .output_share0(d8_t0_26_s0), .output_share1(d8_t0_26_s1));
  reg_module u_reg_t0_27_d8 (.clk(clk), .input_share0(d7_t0_27_s0), .input_share1(d7_t0_27_s1), .output_share0(d8_t0_27_s0), .output_share1(d8_t0_27_s1));
  reg_module u_reg_t0_28_d8 (.clk(clk), .input_share0(d7_t0_28_s0), .input_share1(d7_t0_28_s1), .output_share0(d8_t0_28_s0), .output_share1(d8_t0_28_s1));
  reg_module u_reg_t0_29_d8 (.clk(clk), .input_share0(d7_t0_29_s0), .input_share1(d7_t0_29_s1), .output_share0(d8_t0_29_s0), .output_share1(d8_t0_29_s1));
  reg_module u_reg_t0_30_d8 (.clk(clk), .input_share0(d7_t0_30_s0), .input_share1(d7_t0_30_s1), .output_share0(d8_t0_30_s0), .output_share1(d8_t0_30_s1));
  reg_module u_reg_t0_31_d8 (.clk(clk), .input_share0(d7_t0_31_s0), .input_share1(d7_t0_31_s1), .output_share0(d8_t0_31_s0), .output_share1(d8_t0_31_s1));
  reg_module u_reg_t0_8_d8 (.clk(clk), .input_share0(d7_t0_8_s0), .input_share1(d7_t0_8_s1), .output_share0(d8_t0_8_s0), .output_share1(d8_t0_8_s1));
  reg_module u_reg_t0_9_d8 (.clk(clk), .input_share0(d7_t0_9_s0), .input_share1(d7_t0_9_s1), .output_share0(d8_t0_9_s0), .output_share1(d8_t0_9_s1));
  xor_module u_xor_c8_d8 (.x_share0(d8_i7_s0), .x_share1(d8_i7_s1), .y_share0(d8_t2_7_s0), .y_share1(d8_t2_7_s1), .z_share0(d8_c8_s0), .z_share1(d8_c8_s1));
  xor_module u_xor_o8_d8 (.x_share0(d8_t0_8_s0), .x_share1(d8_t0_8_s1), .y_share0(d8_c8_s0), .y_share1(d8_c8_s1), .z_share0(d8_o8_s0), .z_share1(d8_o8_s1));
  xor_module u_xor_t1_8_d8 (.x_share0(d8_i8_s0), .x_share1(d8_i8_s1), .y_share0(d8_c8_s0), .y_share1(d8_c8_s1), .z_share0(d8_t1_8_s0), .z_share1(d8_t1_8_s1));
  and_module u_and_t2_7_d8 (.clk(clk), .x_share0(d7_t0_7_s0), .x_share1(d7_t0_7_s1), .y_share0(d7_t1_7_s0), .y_share1(d7_t1_7_s1), .rand(r_t2_7), .z_share0(d8_t2_7_s0), .z_share1(d8_t2_7_s1));
  assign r_t2_7 = stage8_share0[2];
  reg_module u_reg_i10_d9 (.clk(clk), .input_share0(d8_i10_s0), .input_share1(d8_i10_s1), .output_share0(d9_i10_s0), .output_share1(d9_i10_s1));
  reg_module u_reg_i11_d9 (.clk(clk), .input_share0(d8_i11_s0), .input_share1(d8_i11_s1), .output_share0(d9_i11_s0), .output_share1(d9_i11_s1));
  reg_module u_reg_i12_d9 (.clk(clk), .input_share0(d8_i12_s0), .input_share1(d8_i12_s1), .output_share0(d9_i12_s0), .output_share1(d9_i12_s1));
  reg_module u_reg_i13_d9 (.clk(clk), .input_share0(d8_i13_s0), .input_share1(d8_i13_s1), .output_share0(d9_i13_s0), .output_share1(d9_i13_s1));
  reg_module u_reg_i14_d9 (.clk(clk), .input_share0(d8_i14_s0), .input_share1(d8_i14_s1), .output_share0(d9_i14_s0), .output_share1(d9_i14_s1));
  reg_module u_reg_i15_d9 (.clk(clk), .input_share0(d8_i15_s0), .input_share1(d8_i15_s1), .output_share0(d9_i15_s0), .output_share1(d9_i15_s1));
  reg_module u_reg_i16_d9 (.clk(clk), .input_share0(d8_i16_s0), .input_share1(d8_i16_s1), .output_share0(d9_i16_s0), .output_share1(d9_i16_s1));
  reg_module u_reg_i17_d9 (.clk(clk), .input_share0(d8_i17_s0), .input_share1(d8_i17_s1), .output_share0(d9_i17_s0), .output_share1(d9_i17_s1));
  reg_module u_reg_i18_d9 (.clk(clk), .input_share0(d8_i18_s0), .input_share1(d8_i18_s1), .output_share0(d9_i18_s0), .output_share1(d9_i18_s1));
  reg_module u_reg_i19_d9 (.clk(clk), .input_share0(d8_i19_s0), .input_share1(d8_i19_s1), .output_share0(d9_i19_s0), .output_share1(d9_i19_s1));
  reg_module u_reg_i20_d9 (.clk(clk), .input_share0(d8_i20_s0), .input_share1(d8_i20_s1), .output_share0(d9_i20_s0), .output_share1(d9_i20_s1));
  reg_module u_reg_i21_d9 (.clk(clk), .input_share0(d8_i21_s0), .input_share1(d8_i21_s1), .output_share0(d9_i21_s0), .output_share1(d9_i21_s1));
  reg_module u_reg_i22_d9 (.clk(clk), .input_share0(d8_i22_s0), .input_share1(d8_i22_s1), .output_share0(d9_i22_s0), .output_share1(d9_i22_s1));
  reg_module u_reg_i23_d9 (.clk(clk), .input_share0(d8_i23_s0), .input_share1(d8_i23_s1), .output_share0(d9_i23_s0), .output_share1(d9_i23_s1));
  reg_module u_reg_i24_d9 (.clk(clk), .input_share0(d8_i24_s0), .input_share1(d8_i24_s1), .output_share0(d9_i24_s0), .output_share1(d9_i24_s1));
  reg_module u_reg_i25_d9 (.clk(clk), .input_share0(d8_i25_s0), .input_share1(d8_i25_s1), .output_share0(d9_i25_s0), .output_share1(d9_i25_s1));
  reg_module u_reg_i26_d9 (.clk(clk), .input_share0(d8_i26_s0), .input_share1(d8_i26_s1), .output_share0(d9_i26_s0), .output_share1(d9_i26_s1));
  reg_module u_reg_i27_d9 (.clk(clk), .input_share0(d8_i27_s0), .input_share1(d8_i27_s1), .output_share0(d9_i27_s0), .output_share1(d9_i27_s1));
  reg_module u_reg_i28_d9 (.clk(clk), .input_share0(d8_i28_s0), .input_share1(d8_i28_s1), .output_share0(d9_i28_s0), .output_share1(d9_i28_s1));
  reg_module u_reg_i29_d9 (.clk(clk), .input_share0(d8_i29_s0), .input_share1(d8_i29_s1), .output_share0(d9_i29_s0), .output_share1(d9_i29_s1));
  reg_module u_reg_i30_d9 (.clk(clk), .input_share0(d8_i30_s0), .input_share1(d8_i30_s1), .output_share0(d9_i30_s0), .output_share1(d9_i30_s1));
  reg_module u_reg_i8_d9 (.clk(clk), .input_share0(d8_i8_s0), .input_share1(d8_i8_s1), .output_share0(d9_i8_s0), .output_share1(d9_i8_s1));
  reg_module u_reg_i9_d9 (.clk(clk), .input_share0(d8_i9_s0), .input_share1(d8_i9_s1), .output_share0(d9_i9_s0), .output_share1(d9_i9_s1));
  reg_module u_reg_t0_10_d9 (.clk(clk), .input_share0(d8_t0_10_s0), .input_share1(d8_t0_10_s1), .output_share0(d9_t0_10_s0), .output_share1(d9_t0_10_s1));
  reg_module u_reg_t0_11_d9 (.clk(clk), .input_share0(d8_t0_11_s0), .input_share1(d8_t0_11_s1), .output_share0(d9_t0_11_s0), .output_share1(d9_t0_11_s1));
  reg_module u_reg_t0_12_d9 (.clk(clk), .input_share0(d8_t0_12_s0), .input_share1(d8_t0_12_s1), .output_share0(d9_t0_12_s0), .output_share1(d9_t0_12_s1));
  reg_module u_reg_t0_13_d9 (.clk(clk), .input_share0(d8_t0_13_s0), .input_share1(d8_t0_13_s1), .output_share0(d9_t0_13_s0), .output_share1(d9_t0_13_s1));
  reg_module u_reg_t0_14_d9 (.clk(clk), .input_share0(d8_t0_14_s0), .input_share1(d8_t0_14_s1), .output_share0(d9_t0_14_s0), .output_share1(d9_t0_14_s1));
  reg_module u_reg_t0_15_d9 (.clk(clk), .input_share0(d8_t0_15_s0), .input_share1(d8_t0_15_s1), .output_share0(d9_t0_15_s0), .output_share1(d9_t0_15_s1));
  reg_module u_reg_t0_16_d9 (.clk(clk), .input_share0(d8_t0_16_s0), .input_share1(d8_t0_16_s1), .output_share0(d9_t0_16_s0), .output_share1(d9_t0_16_s1));
  reg_module u_reg_t0_17_d9 (.clk(clk), .input_share0(d8_t0_17_s0), .input_share1(d8_t0_17_s1), .output_share0(d9_t0_17_s0), .output_share1(d9_t0_17_s1));
  reg_module u_reg_t0_18_d9 (.clk(clk), .input_share0(d8_t0_18_s0), .input_share1(d8_t0_18_s1), .output_share0(d9_t0_18_s0), .output_share1(d9_t0_18_s1));
  reg_module u_reg_t0_19_d9 (.clk(clk), .input_share0(d8_t0_19_s0), .input_share1(d8_t0_19_s1), .output_share0(d9_t0_19_s0), .output_share1(d9_t0_19_s1));
  reg_module u_reg_t0_20_d9 (.clk(clk), .input_share0(d8_t0_20_s0), .input_share1(d8_t0_20_s1), .output_share0(d9_t0_20_s0), .output_share1(d9_t0_20_s1));
  reg_module u_reg_t0_21_d9 (.clk(clk), .input_share0(d8_t0_21_s0), .input_share1(d8_t0_21_s1), .output_share0(d9_t0_21_s0), .output_share1(d9_t0_21_s1));
  reg_module u_reg_t0_22_d9 (.clk(clk), .input_share0(d8_t0_22_s0), .input_share1(d8_t0_22_s1), .output_share0(d9_t0_22_s0), .output_share1(d9_t0_22_s1));
  reg_module u_reg_t0_23_d9 (.clk(clk), .input_share0(d8_t0_23_s0), .input_share1(d8_t0_23_s1), .output_share0(d9_t0_23_s0), .output_share1(d9_t0_23_s1));
  reg_module u_reg_t0_24_d9 (.clk(clk), .input_share0(d8_t0_24_s0), .input_share1(d8_t0_24_s1), .output_share0(d9_t0_24_s0), .output_share1(d9_t0_24_s1));
  reg_module u_reg_t0_25_d9 (.clk(clk), .input_share0(d8_t0_25_s0), .input_share1(d8_t0_25_s1), .output_share0(d9_t0_25_s0), .output_share1(d9_t0_25_s1));
  reg_module u_reg_t0_26_d9 (.clk(clk), .input_share0(d8_t0_26_s0), .input_share1(d8_t0_26_s1), .output_share0(d9_t0_26_s0), .output_share1(d9_t0_26_s1));
  reg_module u_reg_t0_27_d9 (.clk(clk), .input_share0(d8_t0_27_s0), .input_share1(d8_t0_27_s1), .output_share0(d9_t0_27_s0), .output_share1(d9_t0_27_s1));
  reg_module u_reg_t0_28_d9 (.clk(clk), .input_share0(d8_t0_28_s0), .input_share1(d8_t0_28_s1), .output_share0(d9_t0_28_s0), .output_share1(d9_t0_28_s1));
  reg_module u_reg_t0_29_d9 (.clk(clk), .input_share0(d8_t0_29_s0), .input_share1(d8_t0_29_s1), .output_share0(d9_t0_29_s0), .output_share1(d9_t0_29_s1));
  reg_module u_reg_t0_30_d9 (.clk(clk), .input_share0(d8_t0_30_s0), .input_share1(d8_t0_30_s1), .output_share0(d9_t0_30_s0), .output_share1(d9_t0_30_s1));
  reg_module u_reg_t0_31_d9 (.clk(clk), .input_share0(d8_t0_31_s0), .input_share1(d8_t0_31_s1), .output_share0(d9_t0_31_s0), .output_share1(d9_t0_31_s1));
  reg_module u_reg_t0_9_d9 (.clk(clk), .input_share0(d8_t0_9_s0), .input_share1(d8_t0_9_s1), .output_share0(d9_t0_9_s0), .output_share1(d9_t0_9_s1));
  xor_module u_xor_c9_d9 (.x_share0(d9_i8_s0), .x_share1(d9_i8_s1), .y_share0(d9_t2_8_s0), .y_share1(d9_t2_8_s1), .z_share0(d9_c9_s0), .z_share1(d9_c9_s1));
  xor_module u_xor_o9_d9 (.x_share0(d9_t0_9_s0), .x_share1(d9_t0_9_s1), .y_share0(d9_c9_s0), .y_share1(d9_c9_s1), .z_share0(d9_o9_s0), .z_share1(d9_o9_s1));
  xor_module u_xor_t1_9_d9 (.x_share0(d9_i9_s0), .x_share1(d9_i9_s1), .y_share0(d9_c9_s0), .y_share1(d9_c9_s1), .z_share0(d9_t1_9_s0), .z_share1(d9_t1_9_s1));
  and_module u_and_t2_8_d9 (.clk(clk), .x_share0(d8_t0_8_s0), .x_share1(d8_t0_8_s1), .y_share0(d8_t1_8_s0), .y_share1(d8_t1_8_s1), .rand(r_t2_8), .z_share0(d9_t2_8_s0), .z_share1(d9_t2_8_s1));
  assign r_t2_8 = stage9_share0[0];
  reg_module u_reg_i10_d10 (.clk(clk), .input_share0(d9_i10_s0), .input_share1(d9_i10_s1), .output_share0(d10_i10_s0), .output_share1(d10_i10_s1));
  reg_module u_reg_i11_d10 (.clk(clk), .input_share0(d9_i11_s0), .input_share1(d9_i11_s1), .output_share0(d10_i11_s0), .output_share1(d10_i11_s1));
  reg_module u_reg_i12_d10 (.clk(clk), .input_share0(d9_i12_s0), .input_share1(d9_i12_s1), .output_share0(d10_i12_s0), .output_share1(d10_i12_s1));
  reg_module u_reg_i13_d10 (.clk(clk), .input_share0(d9_i13_s0), .input_share1(d9_i13_s1), .output_share0(d10_i13_s0), .output_share1(d10_i13_s1));
  reg_module u_reg_i14_d10 (.clk(clk), .input_share0(d9_i14_s0), .input_share1(d9_i14_s1), .output_share0(d10_i14_s0), .output_share1(d10_i14_s1));
  reg_module u_reg_i15_d10 (.clk(clk), .input_share0(d9_i15_s0), .input_share1(d9_i15_s1), .output_share0(d10_i15_s0), .output_share1(d10_i15_s1));
  reg_module u_reg_i16_d10 (.clk(clk), .input_share0(d9_i16_s0), .input_share1(d9_i16_s1), .output_share0(d10_i16_s0), .output_share1(d10_i16_s1));
  reg_module u_reg_i17_d10 (.clk(clk), .input_share0(d9_i17_s0), .input_share1(d9_i17_s1), .output_share0(d10_i17_s0), .output_share1(d10_i17_s1));
  reg_module u_reg_i18_d10 (.clk(clk), .input_share0(d9_i18_s0), .input_share1(d9_i18_s1), .output_share0(d10_i18_s0), .output_share1(d10_i18_s1));
  reg_module u_reg_i19_d10 (.clk(clk), .input_share0(d9_i19_s0), .input_share1(d9_i19_s1), .output_share0(d10_i19_s0), .output_share1(d10_i19_s1));
  reg_module u_reg_i20_d10 (.clk(clk), .input_share0(d9_i20_s0), .input_share1(d9_i20_s1), .output_share0(d10_i20_s0), .output_share1(d10_i20_s1));
  reg_module u_reg_i21_d10 (.clk(clk), .input_share0(d9_i21_s0), .input_share1(d9_i21_s1), .output_share0(d10_i21_s0), .output_share1(d10_i21_s1));
  reg_module u_reg_i22_d10 (.clk(clk), .input_share0(d9_i22_s0), .input_share1(d9_i22_s1), .output_share0(d10_i22_s0), .output_share1(d10_i22_s1));
  reg_module u_reg_i23_d10 (.clk(clk), .input_share0(d9_i23_s0), .input_share1(d9_i23_s1), .output_share0(d10_i23_s0), .output_share1(d10_i23_s1));
  reg_module u_reg_i24_d10 (.clk(clk), .input_share0(d9_i24_s0), .input_share1(d9_i24_s1), .output_share0(d10_i24_s0), .output_share1(d10_i24_s1));
  reg_module u_reg_i25_d10 (.clk(clk), .input_share0(d9_i25_s0), .input_share1(d9_i25_s1), .output_share0(d10_i25_s0), .output_share1(d10_i25_s1));
  reg_module u_reg_i26_d10 (.clk(clk), .input_share0(d9_i26_s0), .input_share1(d9_i26_s1), .output_share0(d10_i26_s0), .output_share1(d10_i26_s1));
  reg_module u_reg_i27_d10 (.clk(clk), .input_share0(d9_i27_s0), .input_share1(d9_i27_s1), .output_share0(d10_i27_s0), .output_share1(d10_i27_s1));
  reg_module u_reg_i28_d10 (.clk(clk), .input_share0(d9_i28_s0), .input_share1(d9_i28_s1), .output_share0(d10_i28_s0), .output_share1(d10_i28_s1));
  reg_module u_reg_i29_d10 (.clk(clk), .input_share0(d9_i29_s0), .input_share1(d9_i29_s1), .output_share0(d10_i29_s0), .output_share1(d10_i29_s1));
  reg_module u_reg_i30_d10 (.clk(clk), .input_share0(d9_i30_s0), .input_share1(d9_i30_s1), .output_share0(d10_i30_s0), .output_share1(d10_i30_s1));
  reg_module u_reg_i9_d10 (.clk(clk), .input_share0(d9_i9_s0), .input_share1(d9_i9_s1), .output_share0(d10_i9_s0), .output_share1(d10_i9_s1));
  reg_module u_reg_t0_10_d10 (.clk(clk), .input_share0(d9_t0_10_s0), .input_share1(d9_t0_10_s1), .output_share0(d10_t0_10_s0), .output_share1(d10_t0_10_s1));
  reg_module u_reg_t0_11_d10 (.clk(clk), .input_share0(d9_t0_11_s0), .input_share1(d9_t0_11_s1), .output_share0(d10_t0_11_s0), .output_share1(d10_t0_11_s1));
  reg_module u_reg_t0_12_d10 (.clk(clk), .input_share0(d9_t0_12_s0), .input_share1(d9_t0_12_s1), .output_share0(d10_t0_12_s0), .output_share1(d10_t0_12_s1));
  reg_module u_reg_t0_13_d10 (.clk(clk), .input_share0(d9_t0_13_s0), .input_share1(d9_t0_13_s1), .output_share0(d10_t0_13_s0), .output_share1(d10_t0_13_s1));
  reg_module u_reg_t0_14_d10 (.clk(clk), .input_share0(d9_t0_14_s0), .input_share1(d9_t0_14_s1), .output_share0(d10_t0_14_s0), .output_share1(d10_t0_14_s1));
  reg_module u_reg_t0_15_d10 (.clk(clk), .input_share0(d9_t0_15_s0), .input_share1(d9_t0_15_s1), .output_share0(d10_t0_15_s0), .output_share1(d10_t0_15_s1));
  reg_module u_reg_t0_16_d10 (.clk(clk), .input_share0(d9_t0_16_s0), .input_share1(d9_t0_16_s1), .output_share0(d10_t0_16_s0), .output_share1(d10_t0_16_s1));
  reg_module u_reg_t0_17_d10 (.clk(clk), .input_share0(d9_t0_17_s0), .input_share1(d9_t0_17_s1), .output_share0(d10_t0_17_s0), .output_share1(d10_t0_17_s1));
  reg_module u_reg_t0_18_d10 (.clk(clk), .input_share0(d9_t0_18_s0), .input_share1(d9_t0_18_s1), .output_share0(d10_t0_18_s0), .output_share1(d10_t0_18_s1));
  reg_module u_reg_t0_19_d10 (.clk(clk), .input_share0(d9_t0_19_s0), .input_share1(d9_t0_19_s1), .output_share0(d10_t0_19_s0), .output_share1(d10_t0_19_s1));
  reg_module u_reg_t0_20_d10 (.clk(clk), .input_share0(d9_t0_20_s0), .input_share1(d9_t0_20_s1), .output_share0(d10_t0_20_s0), .output_share1(d10_t0_20_s1));
  reg_module u_reg_t0_21_d10 (.clk(clk), .input_share0(d9_t0_21_s0), .input_share1(d9_t0_21_s1), .output_share0(d10_t0_21_s0), .output_share1(d10_t0_21_s1));
  reg_module u_reg_t0_22_d10 (.clk(clk), .input_share0(d9_t0_22_s0), .input_share1(d9_t0_22_s1), .output_share0(d10_t0_22_s0), .output_share1(d10_t0_22_s1));
  reg_module u_reg_t0_23_d10 (.clk(clk), .input_share0(d9_t0_23_s0), .input_share1(d9_t0_23_s1), .output_share0(d10_t0_23_s0), .output_share1(d10_t0_23_s1));
  reg_module u_reg_t0_24_d10 (.clk(clk), .input_share0(d9_t0_24_s0), .input_share1(d9_t0_24_s1), .output_share0(d10_t0_24_s0), .output_share1(d10_t0_24_s1));
  reg_module u_reg_t0_25_d10 (.clk(clk), .input_share0(d9_t0_25_s0), .input_share1(d9_t0_25_s1), .output_share0(d10_t0_25_s0), .output_share1(d10_t0_25_s1));
  reg_module u_reg_t0_26_d10 (.clk(clk), .input_share0(d9_t0_26_s0), .input_share1(d9_t0_26_s1), .output_share0(d10_t0_26_s0), .output_share1(d10_t0_26_s1));
  reg_module u_reg_t0_27_d10 (.clk(clk), .input_share0(d9_t0_27_s0), .input_share1(d9_t0_27_s1), .output_share0(d10_t0_27_s0), .output_share1(d10_t0_27_s1));
  reg_module u_reg_t0_28_d10 (.clk(clk), .input_share0(d9_t0_28_s0), .input_share1(d9_t0_28_s1), .output_share0(d10_t0_28_s0), .output_share1(d10_t0_28_s1));
  reg_module u_reg_t0_29_d10 (.clk(clk), .input_share0(d9_t0_29_s0), .input_share1(d9_t0_29_s1), .output_share0(d10_t0_29_s0), .output_share1(d10_t0_29_s1));
  reg_module u_reg_t0_30_d10 (.clk(clk), .input_share0(d9_t0_30_s0), .input_share1(d9_t0_30_s1), .output_share0(d10_t0_30_s0), .output_share1(d10_t0_30_s1));
  reg_module u_reg_t0_31_d10 (.clk(clk), .input_share0(d9_t0_31_s0), .input_share1(d9_t0_31_s1), .output_share0(d10_t0_31_s0), .output_share1(d10_t0_31_s1));
  xor_module u_xor_c10_d10 (.x_share0(d10_i9_s0), .x_share1(d10_i9_s1), .y_share0(d10_t2_9_s0), .y_share1(d10_t2_9_s1), .z_share0(d10_c10_s0), .z_share1(d10_c10_s1));
  xor_module u_xor_o10_d10 (.x_share0(d10_t0_10_s0), .x_share1(d10_t0_10_s1), .y_share0(d10_c10_s0), .y_share1(d10_c10_s1), .z_share0(d10_o10_s0), .z_share1(d10_o10_s1));
  xor_module u_xor_t1_10_d10 (.x_share0(d10_i10_s0), .x_share1(d10_i10_s1), .y_share0(d10_c10_s0), .y_share1(d10_c10_s1), .z_share0(d10_t1_10_s0), .z_share1(d10_t1_10_s1));
  and_module u_and_t2_9_d10 (.clk(clk), .x_share0(d9_t0_9_s0), .x_share1(d9_t0_9_s1), .y_share0(d9_t1_9_s0), .y_share1(d9_t1_9_s1), .rand(r_t2_9), .z_share0(d10_t2_9_s0), .z_share1(d10_t2_9_s1));
  assign r_t2_9 = stage10_share0[1];
  reg_module u_reg_i10_d11 (.clk(clk), .input_share0(d10_i10_s0), .input_share1(d10_i10_s1), .output_share0(d11_i10_s0), .output_share1(d11_i10_s1));
  reg_module u_reg_i11_d11 (.clk(clk), .input_share0(d10_i11_s0), .input_share1(d10_i11_s1), .output_share0(d11_i11_s0), .output_share1(d11_i11_s1));
  reg_module u_reg_i12_d11 (.clk(clk), .input_share0(d10_i12_s0), .input_share1(d10_i12_s1), .output_share0(d11_i12_s0), .output_share1(d11_i12_s1));
  reg_module u_reg_i13_d11 (.clk(clk), .input_share0(d10_i13_s0), .input_share1(d10_i13_s1), .output_share0(d11_i13_s0), .output_share1(d11_i13_s1));
  reg_module u_reg_i14_d11 (.clk(clk), .input_share0(d10_i14_s0), .input_share1(d10_i14_s1), .output_share0(d11_i14_s0), .output_share1(d11_i14_s1));
  reg_module u_reg_i15_d11 (.clk(clk), .input_share0(d10_i15_s0), .input_share1(d10_i15_s1), .output_share0(d11_i15_s0), .output_share1(d11_i15_s1));
  reg_module u_reg_i16_d11 (.clk(clk), .input_share0(d10_i16_s0), .input_share1(d10_i16_s1), .output_share0(d11_i16_s0), .output_share1(d11_i16_s1));
  reg_module u_reg_i17_d11 (.clk(clk), .input_share0(d10_i17_s0), .input_share1(d10_i17_s1), .output_share0(d11_i17_s0), .output_share1(d11_i17_s1));
  reg_module u_reg_i18_d11 (.clk(clk), .input_share0(d10_i18_s0), .input_share1(d10_i18_s1), .output_share0(d11_i18_s0), .output_share1(d11_i18_s1));
  reg_module u_reg_i19_d11 (.clk(clk), .input_share0(d10_i19_s0), .input_share1(d10_i19_s1), .output_share0(d11_i19_s0), .output_share1(d11_i19_s1));
  reg_module u_reg_i20_d11 (.clk(clk), .input_share0(d10_i20_s0), .input_share1(d10_i20_s1), .output_share0(d11_i20_s0), .output_share1(d11_i20_s1));
  reg_module u_reg_i21_d11 (.clk(clk), .input_share0(d10_i21_s0), .input_share1(d10_i21_s1), .output_share0(d11_i21_s0), .output_share1(d11_i21_s1));
  reg_module u_reg_i22_d11 (.clk(clk), .input_share0(d10_i22_s0), .input_share1(d10_i22_s1), .output_share0(d11_i22_s0), .output_share1(d11_i22_s1));
  reg_module u_reg_i23_d11 (.clk(clk), .input_share0(d10_i23_s0), .input_share1(d10_i23_s1), .output_share0(d11_i23_s0), .output_share1(d11_i23_s1));
  reg_module u_reg_i24_d11 (.clk(clk), .input_share0(d10_i24_s0), .input_share1(d10_i24_s1), .output_share0(d11_i24_s0), .output_share1(d11_i24_s1));
  reg_module u_reg_i25_d11 (.clk(clk), .input_share0(d10_i25_s0), .input_share1(d10_i25_s1), .output_share0(d11_i25_s0), .output_share1(d11_i25_s1));
  reg_module u_reg_i26_d11 (.clk(clk), .input_share0(d10_i26_s0), .input_share1(d10_i26_s1), .output_share0(d11_i26_s0), .output_share1(d11_i26_s1));
  reg_module u_reg_i27_d11 (.clk(clk), .input_share0(d10_i27_s0), .input_share1(d10_i27_s1), .output_share0(d11_i27_s0), .output_share1(d11_i27_s1));
  reg_module u_reg_i28_d11 (.clk(clk), .input_share0(d10_i28_s0), .input_share1(d10_i28_s1), .output_share0(d11_i28_s0), .output_share1(d11_i28_s1));
  reg_module u_reg_i29_d11 (.clk(clk), .input_share0(d10_i29_s0), .input_share1(d10_i29_s1), .output_share0(d11_i29_s0), .output_share1(d11_i29_s1));
  reg_module u_reg_i30_d11 (.clk(clk), .input_share0(d10_i30_s0), .input_share1(d10_i30_s1), .output_share0(d11_i30_s0), .output_share1(d11_i30_s1));
  reg_module u_reg_t0_11_d11 (.clk(clk), .input_share0(d10_t0_11_s0), .input_share1(d10_t0_11_s1), .output_share0(d11_t0_11_s0), .output_share1(d11_t0_11_s1));
  reg_module u_reg_t0_12_d11 (.clk(clk), .input_share0(d10_t0_12_s0), .input_share1(d10_t0_12_s1), .output_share0(d11_t0_12_s0), .output_share1(d11_t0_12_s1));
  reg_module u_reg_t0_13_d11 (.clk(clk), .input_share0(d10_t0_13_s0), .input_share1(d10_t0_13_s1), .output_share0(d11_t0_13_s0), .output_share1(d11_t0_13_s1));
  reg_module u_reg_t0_14_d11 (.clk(clk), .input_share0(d10_t0_14_s0), .input_share1(d10_t0_14_s1), .output_share0(d11_t0_14_s0), .output_share1(d11_t0_14_s1));
  reg_module u_reg_t0_15_d11 (.clk(clk), .input_share0(d10_t0_15_s0), .input_share1(d10_t0_15_s1), .output_share0(d11_t0_15_s0), .output_share1(d11_t0_15_s1));
  reg_module u_reg_t0_16_d11 (.clk(clk), .input_share0(d10_t0_16_s0), .input_share1(d10_t0_16_s1), .output_share0(d11_t0_16_s0), .output_share1(d11_t0_16_s1));
  reg_module u_reg_t0_17_d11 (.clk(clk), .input_share0(d10_t0_17_s0), .input_share1(d10_t0_17_s1), .output_share0(d11_t0_17_s0), .output_share1(d11_t0_17_s1));
  reg_module u_reg_t0_18_d11 (.clk(clk), .input_share0(d10_t0_18_s0), .input_share1(d10_t0_18_s1), .output_share0(d11_t0_18_s0), .output_share1(d11_t0_18_s1));
  reg_module u_reg_t0_19_d11 (.clk(clk), .input_share0(d10_t0_19_s0), .input_share1(d10_t0_19_s1), .output_share0(d11_t0_19_s0), .output_share1(d11_t0_19_s1));
  reg_module u_reg_t0_20_d11 (.clk(clk), .input_share0(d10_t0_20_s0), .input_share1(d10_t0_20_s1), .output_share0(d11_t0_20_s0), .output_share1(d11_t0_20_s1));
  reg_module u_reg_t0_21_d11 (.clk(clk), .input_share0(d10_t0_21_s0), .input_share1(d10_t0_21_s1), .output_share0(d11_t0_21_s0), .output_share1(d11_t0_21_s1));
  reg_module u_reg_t0_22_d11 (.clk(clk), .input_share0(d10_t0_22_s0), .input_share1(d10_t0_22_s1), .output_share0(d11_t0_22_s0), .output_share1(d11_t0_22_s1));
  reg_module u_reg_t0_23_d11 (.clk(clk), .input_share0(d10_t0_23_s0), .input_share1(d10_t0_23_s1), .output_share0(d11_t0_23_s0), .output_share1(d11_t0_23_s1));
  reg_module u_reg_t0_24_d11 (.clk(clk), .input_share0(d10_t0_24_s0), .input_share1(d10_t0_24_s1), .output_share0(d11_t0_24_s0), .output_share1(d11_t0_24_s1));
  reg_module u_reg_t0_25_d11 (.clk(clk), .input_share0(d10_t0_25_s0), .input_share1(d10_t0_25_s1), .output_share0(d11_t0_25_s0), .output_share1(d11_t0_25_s1));
  reg_module u_reg_t0_26_d11 (.clk(clk), .input_share0(d10_t0_26_s0), .input_share1(d10_t0_26_s1), .output_share0(d11_t0_26_s0), .output_share1(d11_t0_26_s1));
  reg_module u_reg_t0_27_d11 (.clk(clk), .input_share0(d10_t0_27_s0), .input_share1(d10_t0_27_s1), .output_share0(d11_t0_27_s0), .output_share1(d11_t0_27_s1));
  reg_module u_reg_t0_28_d11 (.clk(clk), .input_share0(d10_t0_28_s0), .input_share1(d10_t0_28_s1), .output_share0(d11_t0_28_s0), .output_share1(d11_t0_28_s1));
  reg_module u_reg_t0_29_d11 (.clk(clk), .input_share0(d10_t0_29_s0), .input_share1(d10_t0_29_s1), .output_share0(d11_t0_29_s0), .output_share1(d11_t0_29_s1));
  reg_module u_reg_t0_30_d11 (.clk(clk), .input_share0(d10_t0_30_s0), .input_share1(d10_t0_30_s1), .output_share0(d11_t0_30_s0), .output_share1(d11_t0_30_s1));
  reg_module u_reg_t0_31_d11 (.clk(clk), .input_share0(d10_t0_31_s0), .input_share1(d10_t0_31_s1), .output_share0(d11_t0_31_s0), .output_share1(d11_t0_31_s1));
  xor_module u_xor_c11_d11 (.x_share0(d11_i10_s0), .x_share1(d11_i10_s1), .y_share0(d11_t2_10_s0), .y_share1(d11_t2_10_s1), .z_share0(d11_c11_s0), .z_share1(d11_c11_s1));
  xor_module u_xor_o11_d11 (.x_share0(d11_t0_11_s0), .x_share1(d11_t0_11_s1), .y_share0(d11_c11_s0), .y_share1(d11_c11_s1), .z_share0(d11_o11_s0), .z_share1(d11_o11_s1));
  xor_module u_xor_t1_11_d11 (.x_share0(d11_i11_s0), .x_share1(d11_i11_s1), .y_share0(d11_c11_s0), .y_share1(d11_c11_s1), .z_share0(d11_t1_11_s0), .z_share1(d11_t1_11_s1));
  and_module u_and_t2_10_d11 (.clk(clk), .x_share0(d10_t0_10_s0), .x_share1(d10_t0_10_s1), .y_share0(d10_t1_10_s0), .y_share1(d10_t1_10_s1), .rand(r_t2_10), .z_share0(d11_t2_10_s0), .z_share1(d11_t2_10_s1));
  assign r_t2_10 = stage11_share0[2];
  reg_module u_reg_i11_d12 (.clk(clk), .input_share0(d11_i11_s0), .input_share1(d11_i11_s1), .output_share0(d12_i11_s0), .output_share1(d12_i11_s1));
  reg_module u_reg_i12_d12 (.clk(clk), .input_share0(d11_i12_s0), .input_share1(d11_i12_s1), .output_share0(d12_i12_s0), .output_share1(d12_i12_s1));
  reg_module u_reg_i13_d12 (.clk(clk), .input_share0(d11_i13_s0), .input_share1(d11_i13_s1), .output_share0(d12_i13_s0), .output_share1(d12_i13_s1));
  reg_module u_reg_i14_d12 (.clk(clk), .input_share0(d11_i14_s0), .input_share1(d11_i14_s1), .output_share0(d12_i14_s0), .output_share1(d12_i14_s1));
  reg_module u_reg_i15_d12 (.clk(clk), .input_share0(d11_i15_s0), .input_share1(d11_i15_s1), .output_share0(d12_i15_s0), .output_share1(d12_i15_s1));
  reg_module u_reg_i16_d12 (.clk(clk), .input_share0(d11_i16_s0), .input_share1(d11_i16_s1), .output_share0(d12_i16_s0), .output_share1(d12_i16_s1));
  reg_module u_reg_i17_d12 (.clk(clk), .input_share0(d11_i17_s0), .input_share1(d11_i17_s1), .output_share0(d12_i17_s0), .output_share1(d12_i17_s1));
  reg_module u_reg_i18_d12 (.clk(clk), .input_share0(d11_i18_s0), .input_share1(d11_i18_s1), .output_share0(d12_i18_s0), .output_share1(d12_i18_s1));
  reg_module u_reg_i19_d12 (.clk(clk), .input_share0(d11_i19_s0), .input_share1(d11_i19_s1), .output_share0(d12_i19_s0), .output_share1(d12_i19_s1));
  reg_module u_reg_i20_d12 (.clk(clk), .input_share0(d11_i20_s0), .input_share1(d11_i20_s1), .output_share0(d12_i20_s0), .output_share1(d12_i20_s1));
  reg_module u_reg_i21_d12 (.clk(clk), .input_share0(d11_i21_s0), .input_share1(d11_i21_s1), .output_share0(d12_i21_s0), .output_share1(d12_i21_s1));
  reg_module u_reg_i22_d12 (.clk(clk), .input_share0(d11_i22_s0), .input_share1(d11_i22_s1), .output_share0(d12_i22_s0), .output_share1(d12_i22_s1));
  reg_module u_reg_i23_d12 (.clk(clk), .input_share0(d11_i23_s0), .input_share1(d11_i23_s1), .output_share0(d12_i23_s0), .output_share1(d12_i23_s1));
  reg_module u_reg_i24_d12 (.clk(clk), .input_share0(d11_i24_s0), .input_share1(d11_i24_s1), .output_share0(d12_i24_s0), .output_share1(d12_i24_s1));
  reg_module u_reg_i25_d12 (.clk(clk), .input_share0(d11_i25_s0), .input_share1(d11_i25_s1), .output_share0(d12_i25_s0), .output_share1(d12_i25_s1));
  reg_module u_reg_i26_d12 (.clk(clk), .input_share0(d11_i26_s0), .input_share1(d11_i26_s1), .output_share0(d12_i26_s0), .output_share1(d12_i26_s1));
  reg_module u_reg_i27_d12 (.clk(clk), .input_share0(d11_i27_s0), .input_share1(d11_i27_s1), .output_share0(d12_i27_s0), .output_share1(d12_i27_s1));
  reg_module u_reg_i28_d12 (.clk(clk), .input_share0(d11_i28_s0), .input_share1(d11_i28_s1), .output_share0(d12_i28_s0), .output_share1(d12_i28_s1));
  reg_module u_reg_i29_d12 (.clk(clk), .input_share0(d11_i29_s0), .input_share1(d11_i29_s1), .output_share0(d12_i29_s0), .output_share1(d12_i29_s1));
  reg_module u_reg_i30_d12 (.clk(clk), .input_share0(d11_i30_s0), .input_share1(d11_i30_s1), .output_share0(d12_i30_s0), .output_share1(d12_i30_s1));
  reg_module u_reg_t0_12_d12 (.clk(clk), .input_share0(d11_t0_12_s0), .input_share1(d11_t0_12_s1), .output_share0(d12_t0_12_s0), .output_share1(d12_t0_12_s1));
  reg_module u_reg_t0_13_d12 (.clk(clk), .input_share0(d11_t0_13_s0), .input_share1(d11_t0_13_s1), .output_share0(d12_t0_13_s0), .output_share1(d12_t0_13_s1));
  reg_module u_reg_t0_14_d12 (.clk(clk), .input_share0(d11_t0_14_s0), .input_share1(d11_t0_14_s1), .output_share0(d12_t0_14_s0), .output_share1(d12_t0_14_s1));
  reg_module u_reg_t0_15_d12 (.clk(clk), .input_share0(d11_t0_15_s0), .input_share1(d11_t0_15_s1), .output_share0(d12_t0_15_s0), .output_share1(d12_t0_15_s1));
  reg_module u_reg_t0_16_d12 (.clk(clk), .input_share0(d11_t0_16_s0), .input_share1(d11_t0_16_s1), .output_share0(d12_t0_16_s0), .output_share1(d12_t0_16_s1));
  reg_module u_reg_t0_17_d12 (.clk(clk), .input_share0(d11_t0_17_s0), .input_share1(d11_t0_17_s1), .output_share0(d12_t0_17_s0), .output_share1(d12_t0_17_s1));
  reg_module u_reg_t0_18_d12 (.clk(clk), .input_share0(d11_t0_18_s0), .input_share1(d11_t0_18_s1), .output_share0(d12_t0_18_s0), .output_share1(d12_t0_18_s1));
  reg_module u_reg_t0_19_d12 (.clk(clk), .input_share0(d11_t0_19_s0), .input_share1(d11_t0_19_s1), .output_share0(d12_t0_19_s0), .output_share1(d12_t0_19_s1));
  reg_module u_reg_t0_20_d12 (.clk(clk), .input_share0(d11_t0_20_s0), .input_share1(d11_t0_20_s1), .output_share0(d12_t0_20_s0), .output_share1(d12_t0_20_s1));
  reg_module u_reg_t0_21_d12 (.clk(clk), .input_share0(d11_t0_21_s0), .input_share1(d11_t0_21_s1), .output_share0(d12_t0_21_s0), .output_share1(d12_t0_21_s1));
  reg_module u_reg_t0_22_d12 (.clk(clk), .input_share0(d11_t0_22_s0), .input_share1(d11_t0_22_s1), .output_share0(d12_t0_22_s0), .output_share1(d12_t0_22_s1));
  reg_module u_reg_t0_23_d12 (.clk(clk), .input_share0(d11_t0_23_s0), .input_share1(d11_t0_23_s1), .output_share0(d12_t0_23_s0), .output_share1(d12_t0_23_s1));
  reg_module u_reg_t0_24_d12 (.clk(clk), .input_share0(d11_t0_24_s0), .input_share1(d11_t0_24_s1), .output_share0(d12_t0_24_s0), .output_share1(d12_t0_24_s1));
  reg_module u_reg_t0_25_d12 (.clk(clk), .input_share0(d11_t0_25_s0), .input_share1(d11_t0_25_s1), .output_share0(d12_t0_25_s0), .output_share1(d12_t0_25_s1));
  reg_module u_reg_t0_26_d12 (.clk(clk), .input_share0(d11_t0_26_s0), .input_share1(d11_t0_26_s1), .output_share0(d12_t0_26_s0), .output_share1(d12_t0_26_s1));
  reg_module u_reg_t0_27_d12 (.clk(clk), .input_share0(d11_t0_27_s0), .input_share1(d11_t0_27_s1), .output_share0(d12_t0_27_s0), .output_share1(d12_t0_27_s1));
  reg_module u_reg_t0_28_d12 (.clk(clk), .input_share0(d11_t0_28_s0), .input_share1(d11_t0_28_s1), .output_share0(d12_t0_28_s0), .output_share1(d12_t0_28_s1));
  reg_module u_reg_t0_29_d12 (.clk(clk), .input_share0(d11_t0_29_s0), .input_share1(d11_t0_29_s1), .output_share0(d12_t0_29_s0), .output_share1(d12_t0_29_s1));
  reg_module u_reg_t0_30_d12 (.clk(clk), .input_share0(d11_t0_30_s0), .input_share1(d11_t0_30_s1), .output_share0(d12_t0_30_s0), .output_share1(d12_t0_30_s1));
  reg_module u_reg_t0_31_d12 (.clk(clk), .input_share0(d11_t0_31_s0), .input_share1(d11_t0_31_s1), .output_share0(d12_t0_31_s0), .output_share1(d12_t0_31_s1));
  xor_module u_xor_c12_d12 (.x_share0(d12_i11_s0), .x_share1(d12_i11_s1), .y_share0(d12_t2_11_s0), .y_share1(d12_t2_11_s1), .z_share0(d12_c12_s0), .z_share1(d12_c12_s1));
  xor_module u_xor_o12_d12 (.x_share0(d12_t0_12_s0), .x_share1(d12_t0_12_s1), .y_share0(d12_c12_s0), .y_share1(d12_c12_s1), .z_share0(d12_o12_s0), .z_share1(d12_o12_s1));
  xor_module u_xor_t1_12_d12 (.x_share0(d12_i12_s0), .x_share1(d12_i12_s1), .y_share0(d12_c12_s0), .y_share1(d12_c12_s1), .z_share0(d12_t1_12_s0), .z_share1(d12_t1_12_s1));
  and_module u_and_t2_11_d12 (.clk(clk), .x_share0(d11_t0_11_s0), .x_share1(d11_t0_11_s1), .y_share0(d11_t1_11_s0), .y_share1(d11_t1_11_s1), .rand(r_t2_11), .z_share0(d12_t2_11_s0), .z_share1(d12_t2_11_s1));
  assign r_t2_11 = stage12_share0[0];
  reg_module u_reg_i12_d13 (.clk(clk), .input_share0(d12_i12_s0), .input_share1(d12_i12_s1), .output_share0(d13_i12_s0), .output_share1(d13_i12_s1));
  reg_module u_reg_i13_d13 (.clk(clk), .input_share0(d12_i13_s0), .input_share1(d12_i13_s1), .output_share0(d13_i13_s0), .output_share1(d13_i13_s1));
  reg_module u_reg_i14_d13 (.clk(clk), .input_share0(d12_i14_s0), .input_share1(d12_i14_s1), .output_share0(d13_i14_s0), .output_share1(d13_i14_s1));
  reg_module u_reg_i15_d13 (.clk(clk), .input_share0(d12_i15_s0), .input_share1(d12_i15_s1), .output_share0(d13_i15_s0), .output_share1(d13_i15_s1));
  reg_module u_reg_i16_d13 (.clk(clk), .input_share0(d12_i16_s0), .input_share1(d12_i16_s1), .output_share0(d13_i16_s0), .output_share1(d13_i16_s1));
  reg_module u_reg_i17_d13 (.clk(clk), .input_share0(d12_i17_s0), .input_share1(d12_i17_s1), .output_share0(d13_i17_s0), .output_share1(d13_i17_s1));
  reg_module u_reg_i18_d13 (.clk(clk), .input_share0(d12_i18_s0), .input_share1(d12_i18_s1), .output_share0(d13_i18_s0), .output_share1(d13_i18_s1));
  reg_module u_reg_i19_d13 (.clk(clk), .input_share0(d12_i19_s0), .input_share1(d12_i19_s1), .output_share0(d13_i19_s0), .output_share1(d13_i19_s1));
  reg_module u_reg_i20_d13 (.clk(clk), .input_share0(d12_i20_s0), .input_share1(d12_i20_s1), .output_share0(d13_i20_s0), .output_share1(d13_i20_s1));
  reg_module u_reg_i21_d13 (.clk(clk), .input_share0(d12_i21_s0), .input_share1(d12_i21_s1), .output_share0(d13_i21_s0), .output_share1(d13_i21_s1));
  reg_module u_reg_i22_d13 (.clk(clk), .input_share0(d12_i22_s0), .input_share1(d12_i22_s1), .output_share0(d13_i22_s0), .output_share1(d13_i22_s1));
  reg_module u_reg_i23_d13 (.clk(clk), .input_share0(d12_i23_s0), .input_share1(d12_i23_s1), .output_share0(d13_i23_s0), .output_share1(d13_i23_s1));
  reg_module u_reg_i24_d13 (.clk(clk), .input_share0(d12_i24_s0), .input_share1(d12_i24_s1), .output_share0(d13_i24_s0), .output_share1(d13_i24_s1));
  reg_module u_reg_i25_d13 (.clk(clk), .input_share0(d12_i25_s0), .input_share1(d12_i25_s1), .output_share0(d13_i25_s0), .output_share1(d13_i25_s1));
  reg_module u_reg_i26_d13 (.clk(clk), .input_share0(d12_i26_s0), .input_share1(d12_i26_s1), .output_share0(d13_i26_s0), .output_share1(d13_i26_s1));
  reg_module u_reg_i27_d13 (.clk(clk), .input_share0(d12_i27_s0), .input_share1(d12_i27_s1), .output_share0(d13_i27_s0), .output_share1(d13_i27_s1));
  reg_module u_reg_i28_d13 (.clk(clk), .input_share0(d12_i28_s0), .input_share1(d12_i28_s1), .output_share0(d13_i28_s0), .output_share1(d13_i28_s1));
  reg_module u_reg_i29_d13 (.clk(clk), .input_share0(d12_i29_s0), .input_share1(d12_i29_s1), .output_share0(d13_i29_s0), .output_share1(d13_i29_s1));
  reg_module u_reg_i30_d13 (.clk(clk), .input_share0(d12_i30_s0), .input_share1(d12_i30_s1), .output_share0(d13_i30_s0), .output_share1(d13_i30_s1));
  reg_module u_reg_t0_13_d13 (.clk(clk), .input_share0(d12_t0_13_s0), .input_share1(d12_t0_13_s1), .output_share0(d13_t0_13_s0), .output_share1(d13_t0_13_s1));
  reg_module u_reg_t0_14_d13 (.clk(clk), .input_share0(d12_t0_14_s0), .input_share1(d12_t0_14_s1), .output_share0(d13_t0_14_s0), .output_share1(d13_t0_14_s1));
  reg_module u_reg_t0_15_d13 (.clk(clk), .input_share0(d12_t0_15_s0), .input_share1(d12_t0_15_s1), .output_share0(d13_t0_15_s0), .output_share1(d13_t0_15_s1));
  reg_module u_reg_t0_16_d13 (.clk(clk), .input_share0(d12_t0_16_s0), .input_share1(d12_t0_16_s1), .output_share0(d13_t0_16_s0), .output_share1(d13_t0_16_s1));
  reg_module u_reg_t0_17_d13 (.clk(clk), .input_share0(d12_t0_17_s0), .input_share1(d12_t0_17_s1), .output_share0(d13_t0_17_s0), .output_share1(d13_t0_17_s1));
  reg_module u_reg_t0_18_d13 (.clk(clk), .input_share0(d12_t0_18_s0), .input_share1(d12_t0_18_s1), .output_share0(d13_t0_18_s0), .output_share1(d13_t0_18_s1));
  reg_module u_reg_t0_19_d13 (.clk(clk), .input_share0(d12_t0_19_s0), .input_share1(d12_t0_19_s1), .output_share0(d13_t0_19_s0), .output_share1(d13_t0_19_s1));
  reg_module u_reg_t0_20_d13 (.clk(clk), .input_share0(d12_t0_20_s0), .input_share1(d12_t0_20_s1), .output_share0(d13_t0_20_s0), .output_share1(d13_t0_20_s1));
  reg_module u_reg_t0_21_d13 (.clk(clk), .input_share0(d12_t0_21_s0), .input_share1(d12_t0_21_s1), .output_share0(d13_t0_21_s0), .output_share1(d13_t0_21_s1));
  reg_module u_reg_t0_22_d13 (.clk(clk), .input_share0(d12_t0_22_s0), .input_share1(d12_t0_22_s1), .output_share0(d13_t0_22_s0), .output_share1(d13_t0_22_s1));
  reg_module u_reg_t0_23_d13 (.clk(clk), .input_share0(d12_t0_23_s0), .input_share1(d12_t0_23_s1), .output_share0(d13_t0_23_s0), .output_share1(d13_t0_23_s1));
  reg_module u_reg_t0_24_d13 (.clk(clk), .input_share0(d12_t0_24_s0), .input_share1(d12_t0_24_s1), .output_share0(d13_t0_24_s0), .output_share1(d13_t0_24_s1));
  reg_module u_reg_t0_25_d13 (.clk(clk), .input_share0(d12_t0_25_s0), .input_share1(d12_t0_25_s1), .output_share0(d13_t0_25_s0), .output_share1(d13_t0_25_s1));
  reg_module u_reg_t0_26_d13 (.clk(clk), .input_share0(d12_t0_26_s0), .input_share1(d12_t0_26_s1), .output_share0(d13_t0_26_s0), .output_share1(d13_t0_26_s1));
  reg_module u_reg_t0_27_d13 (.clk(clk), .input_share0(d12_t0_27_s0), .input_share1(d12_t0_27_s1), .output_share0(d13_t0_27_s0), .output_share1(d13_t0_27_s1));
  reg_module u_reg_t0_28_d13 (.clk(clk), .input_share0(d12_t0_28_s0), .input_share1(d12_t0_28_s1), .output_share0(d13_t0_28_s0), .output_share1(d13_t0_28_s1));
  reg_module u_reg_t0_29_d13 (.clk(clk), .input_share0(d12_t0_29_s0), .input_share1(d12_t0_29_s1), .output_share0(d13_t0_29_s0), .output_share1(d13_t0_29_s1));
  reg_module u_reg_t0_30_d13 (.clk(clk), .input_share0(d12_t0_30_s0), .input_share1(d12_t0_30_s1), .output_share0(d13_t0_30_s0), .output_share1(d13_t0_30_s1));
  reg_module u_reg_t0_31_d13 (.clk(clk), .input_share0(d12_t0_31_s0), .input_share1(d12_t0_31_s1), .output_share0(d13_t0_31_s0), .output_share1(d13_t0_31_s1));
  xor_module u_xor_c13_d13 (.x_share0(d13_i12_s0), .x_share1(d13_i12_s1), .y_share0(d13_t2_12_s0), .y_share1(d13_t2_12_s1), .z_share0(d13_c13_s0), .z_share1(d13_c13_s1));
  xor_module u_xor_o13_d13 (.x_share0(d13_t0_13_s0), .x_share1(d13_t0_13_s1), .y_share0(d13_c13_s0), .y_share1(d13_c13_s1), .z_share0(d13_o13_s0), .z_share1(d13_o13_s1));
  xor_module u_xor_t1_13_d13 (.x_share0(d13_i13_s0), .x_share1(d13_i13_s1), .y_share0(d13_c13_s0), .y_share1(d13_c13_s1), .z_share0(d13_t1_13_s0), .z_share1(d13_t1_13_s1));
  and_module u_and_t2_12_d13 (.clk(clk), .x_share0(d12_t0_12_s0), .x_share1(d12_t0_12_s1), .y_share0(d12_t1_12_s0), .y_share1(d12_t1_12_s1), .rand(r_t2_12), .z_share0(d13_t2_12_s0), .z_share1(d13_t2_12_s1));
  assign r_t2_12 = stage13_share0[1];
  reg_module u_reg_i13_d14 (.clk(clk), .input_share0(d13_i13_s0), .input_share1(d13_i13_s1), .output_share0(d14_i13_s0), .output_share1(d14_i13_s1));
  reg_module u_reg_i14_d14 (.clk(clk), .input_share0(d13_i14_s0), .input_share1(d13_i14_s1), .output_share0(d14_i14_s0), .output_share1(d14_i14_s1));
  reg_module u_reg_i15_d14 (.clk(clk), .input_share0(d13_i15_s0), .input_share1(d13_i15_s1), .output_share0(d14_i15_s0), .output_share1(d14_i15_s1));
  reg_module u_reg_i16_d14 (.clk(clk), .input_share0(d13_i16_s0), .input_share1(d13_i16_s1), .output_share0(d14_i16_s0), .output_share1(d14_i16_s1));
  reg_module u_reg_i17_d14 (.clk(clk), .input_share0(d13_i17_s0), .input_share1(d13_i17_s1), .output_share0(d14_i17_s0), .output_share1(d14_i17_s1));
  reg_module u_reg_i18_d14 (.clk(clk), .input_share0(d13_i18_s0), .input_share1(d13_i18_s1), .output_share0(d14_i18_s0), .output_share1(d14_i18_s1));
  reg_module u_reg_i19_d14 (.clk(clk), .input_share0(d13_i19_s0), .input_share1(d13_i19_s1), .output_share0(d14_i19_s0), .output_share1(d14_i19_s1));
  reg_module u_reg_i20_d14 (.clk(clk), .input_share0(d13_i20_s0), .input_share1(d13_i20_s1), .output_share0(d14_i20_s0), .output_share1(d14_i20_s1));
  reg_module u_reg_i21_d14 (.clk(clk), .input_share0(d13_i21_s0), .input_share1(d13_i21_s1), .output_share0(d14_i21_s0), .output_share1(d14_i21_s1));
  reg_module u_reg_i22_d14 (.clk(clk), .input_share0(d13_i22_s0), .input_share1(d13_i22_s1), .output_share0(d14_i22_s0), .output_share1(d14_i22_s1));
  reg_module u_reg_i23_d14 (.clk(clk), .input_share0(d13_i23_s0), .input_share1(d13_i23_s1), .output_share0(d14_i23_s0), .output_share1(d14_i23_s1));
  reg_module u_reg_i24_d14 (.clk(clk), .input_share0(d13_i24_s0), .input_share1(d13_i24_s1), .output_share0(d14_i24_s0), .output_share1(d14_i24_s1));
  reg_module u_reg_i25_d14 (.clk(clk), .input_share0(d13_i25_s0), .input_share1(d13_i25_s1), .output_share0(d14_i25_s0), .output_share1(d14_i25_s1));
  reg_module u_reg_i26_d14 (.clk(clk), .input_share0(d13_i26_s0), .input_share1(d13_i26_s1), .output_share0(d14_i26_s0), .output_share1(d14_i26_s1));
  reg_module u_reg_i27_d14 (.clk(clk), .input_share0(d13_i27_s0), .input_share1(d13_i27_s1), .output_share0(d14_i27_s0), .output_share1(d14_i27_s1));
  reg_module u_reg_i28_d14 (.clk(clk), .input_share0(d13_i28_s0), .input_share1(d13_i28_s1), .output_share0(d14_i28_s0), .output_share1(d14_i28_s1));
  reg_module u_reg_i29_d14 (.clk(clk), .input_share0(d13_i29_s0), .input_share1(d13_i29_s1), .output_share0(d14_i29_s0), .output_share1(d14_i29_s1));
  reg_module u_reg_i30_d14 (.clk(clk), .input_share0(d13_i30_s0), .input_share1(d13_i30_s1), .output_share0(d14_i30_s0), .output_share1(d14_i30_s1));
  reg_module u_reg_t0_14_d14 (.clk(clk), .input_share0(d13_t0_14_s0), .input_share1(d13_t0_14_s1), .output_share0(d14_t0_14_s0), .output_share1(d14_t0_14_s1));
  reg_module u_reg_t0_15_d14 (.clk(clk), .input_share0(d13_t0_15_s0), .input_share1(d13_t0_15_s1), .output_share0(d14_t0_15_s0), .output_share1(d14_t0_15_s1));
  reg_module u_reg_t0_16_d14 (.clk(clk), .input_share0(d13_t0_16_s0), .input_share1(d13_t0_16_s1), .output_share0(d14_t0_16_s0), .output_share1(d14_t0_16_s1));
  reg_module u_reg_t0_17_d14 (.clk(clk), .input_share0(d13_t0_17_s0), .input_share1(d13_t0_17_s1), .output_share0(d14_t0_17_s0), .output_share1(d14_t0_17_s1));
  reg_module u_reg_t0_18_d14 (.clk(clk), .input_share0(d13_t0_18_s0), .input_share1(d13_t0_18_s1), .output_share0(d14_t0_18_s0), .output_share1(d14_t0_18_s1));
  reg_module u_reg_t0_19_d14 (.clk(clk), .input_share0(d13_t0_19_s0), .input_share1(d13_t0_19_s1), .output_share0(d14_t0_19_s0), .output_share1(d14_t0_19_s1));
  reg_module u_reg_t0_20_d14 (.clk(clk), .input_share0(d13_t0_20_s0), .input_share1(d13_t0_20_s1), .output_share0(d14_t0_20_s0), .output_share1(d14_t0_20_s1));
  reg_module u_reg_t0_21_d14 (.clk(clk), .input_share0(d13_t0_21_s0), .input_share1(d13_t0_21_s1), .output_share0(d14_t0_21_s0), .output_share1(d14_t0_21_s1));
  reg_module u_reg_t0_22_d14 (.clk(clk), .input_share0(d13_t0_22_s0), .input_share1(d13_t0_22_s1), .output_share0(d14_t0_22_s0), .output_share1(d14_t0_22_s1));
  reg_module u_reg_t0_23_d14 (.clk(clk), .input_share0(d13_t0_23_s0), .input_share1(d13_t0_23_s1), .output_share0(d14_t0_23_s0), .output_share1(d14_t0_23_s1));
  reg_module u_reg_t0_24_d14 (.clk(clk), .input_share0(d13_t0_24_s0), .input_share1(d13_t0_24_s1), .output_share0(d14_t0_24_s0), .output_share1(d14_t0_24_s1));
  reg_module u_reg_t0_25_d14 (.clk(clk), .input_share0(d13_t0_25_s0), .input_share1(d13_t0_25_s1), .output_share0(d14_t0_25_s0), .output_share1(d14_t0_25_s1));
  reg_module u_reg_t0_26_d14 (.clk(clk), .input_share0(d13_t0_26_s0), .input_share1(d13_t0_26_s1), .output_share0(d14_t0_26_s0), .output_share1(d14_t0_26_s1));
  reg_module u_reg_t0_27_d14 (.clk(clk), .input_share0(d13_t0_27_s0), .input_share1(d13_t0_27_s1), .output_share0(d14_t0_27_s0), .output_share1(d14_t0_27_s1));
  reg_module u_reg_t0_28_d14 (.clk(clk), .input_share0(d13_t0_28_s0), .input_share1(d13_t0_28_s1), .output_share0(d14_t0_28_s0), .output_share1(d14_t0_28_s1));
  reg_module u_reg_t0_29_d14 (.clk(clk), .input_share0(d13_t0_29_s0), .input_share1(d13_t0_29_s1), .output_share0(d14_t0_29_s0), .output_share1(d14_t0_29_s1));
  reg_module u_reg_t0_30_d14 (.clk(clk), .input_share0(d13_t0_30_s0), .input_share1(d13_t0_30_s1), .output_share0(d14_t0_30_s0), .output_share1(d14_t0_30_s1));
  reg_module u_reg_t0_31_d14 (.clk(clk), .input_share0(d13_t0_31_s0), .input_share1(d13_t0_31_s1), .output_share0(d14_t0_31_s0), .output_share1(d14_t0_31_s1));
  xor_module u_xor_c14_d14 (.x_share0(d14_i13_s0), .x_share1(d14_i13_s1), .y_share0(d14_t2_13_s0), .y_share1(d14_t2_13_s1), .z_share0(d14_c14_s0), .z_share1(d14_c14_s1));
  xor_module u_xor_o14_d14 (.x_share0(d14_t0_14_s0), .x_share1(d14_t0_14_s1), .y_share0(d14_c14_s0), .y_share1(d14_c14_s1), .z_share0(d14_o14_s0), .z_share1(d14_o14_s1));
  xor_module u_xor_t1_14_d14 (.x_share0(d14_i14_s0), .x_share1(d14_i14_s1), .y_share0(d14_c14_s0), .y_share1(d14_c14_s1), .z_share0(d14_t1_14_s0), .z_share1(d14_t1_14_s1));
  and_module u_and_t2_13_d14 (.clk(clk), .x_share0(d13_t0_13_s0), .x_share1(d13_t0_13_s1), .y_share0(d13_t1_13_s0), .y_share1(d13_t1_13_s1), .rand(r_t2_13), .z_share0(d14_t2_13_s0), .z_share1(d14_t2_13_s1));
  assign r_t2_13 = stage14_share0[2];
  reg_module u_reg_i14_d15 (.clk(clk), .input_share0(d14_i14_s0), .input_share1(d14_i14_s1), .output_share0(d15_i14_s0), .output_share1(d15_i14_s1));
  reg_module u_reg_i15_d15 (.clk(clk), .input_share0(d14_i15_s0), .input_share1(d14_i15_s1), .output_share0(d15_i15_s0), .output_share1(d15_i15_s1));
  reg_module u_reg_i16_d15 (.clk(clk), .input_share0(d14_i16_s0), .input_share1(d14_i16_s1), .output_share0(d15_i16_s0), .output_share1(d15_i16_s1));
  reg_module u_reg_i17_d15 (.clk(clk), .input_share0(d14_i17_s0), .input_share1(d14_i17_s1), .output_share0(d15_i17_s0), .output_share1(d15_i17_s1));
  reg_module u_reg_i18_d15 (.clk(clk), .input_share0(d14_i18_s0), .input_share1(d14_i18_s1), .output_share0(d15_i18_s0), .output_share1(d15_i18_s1));
  reg_module u_reg_i19_d15 (.clk(clk), .input_share0(d14_i19_s0), .input_share1(d14_i19_s1), .output_share0(d15_i19_s0), .output_share1(d15_i19_s1));
  reg_module u_reg_i20_d15 (.clk(clk), .input_share0(d14_i20_s0), .input_share1(d14_i20_s1), .output_share0(d15_i20_s0), .output_share1(d15_i20_s1));
  reg_module u_reg_i21_d15 (.clk(clk), .input_share0(d14_i21_s0), .input_share1(d14_i21_s1), .output_share0(d15_i21_s0), .output_share1(d15_i21_s1));
  reg_module u_reg_i22_d15 (.clk(clk), .input_share0(d14_i22_s0), .input_share1(d14_i22_s1), .output_share0(d15_i22_s0), .output_share1(d15_i22_s1));
  reg_module u_reg_i23_d15 (.clk(clk), .input_share0(d14_i23_s0), .input_share1(d14_i23_s1), .output_share0(d15_i23_s0), .output_share1(d15_i23_s1));
  reg_module u_reg_i24_d15 (.clk(clk), .input_share0(d14_i24_s0), .input_share1(d14_i24_s1), .output_share0(d15_i24_s0), .output_share1(d15_i24_s1));
  reg_module u_reg_i25_d15 (.clk(clk), .input_share0(d14_i25_s0), .input_share1(d14_i25_s1), .output_share0(d15_i25_s0), .output_share1(d15_i25_s1));
  reg_module u_reg_i26_d15 (.clk(clk), .input_share0(d14_i26_s0), .input_share1(d14_i26_s1), .output_share0(d15_i26_s0), .output_share1(d15_i26_s1));
  reg_module u_reg_i27_d15 (.clk(clk), .input_share0(d14_i27_s0), .input_share1(d14_i27_s1), .output_share0(d15_i27_s0), .output_share1(d15_i27_s1));
  reg_module u_reg_i28_d15 (.clk(clk), .input_share0(d14_i28_s0), .input_share1(d14_i28_s1), .output_share0(d15_i28_s0), .output_share1(d15_i28_s1));
  reg_module u_reg_i29_d15 (.clk(clk), .input_share0(d14_i29_s0), .input_share1(d14_i29_s1), .output_share0(d15_i29_s0), .output_share1(d15_i29_s1));
  reg_module u_reg_i30_d15 (.clk(clk), .input_share0(d14_i30_s0), .input_share1(d14_i30_s1), .output_share0(d15_i30_s0), .output_share1(d15_i30_s1));
  reg_module u_reg_t0_15_d15 (.clk(clk), .input_share0(d14_t0_15_s0), .input_share1(d14_t0_15_s1), .output_share0(d15_t0_15_s0), .output_share1(d15_t0_15_s1));
  reg_module u_reg_t0_16_d15 (.clk(clk), .input_share0(d14_t0_16_s0), .input_share1(d14_t0_16_s1), .output_share0(d15_t0_16_s0), .output_share1(d15_t0_16_s1));
  reg_module u_reg_t0_17_d15 (.clk(clk), .input_share0(d14_t0_17_s0), .input_share1(d14_t0_17_s1), .output_share0(d15_t0_17_s0), .output_share1(d15_t0_17_s1));
  reg_module u_reg_t0_18_d15 (.clk(clk), .input_share0(d14_t0_18_s0), .input_share1(d14_t0_18_s1), .output_share0(d15_t0_18_s0), .output_share1(d15_t0_18_s1));
  reg_module u_reg_t0_19_d15 (.clk(clk), .input_share0(d14_t0_19_s0), .input_share1(d14_t0_19_s1), .output_share0(d15_t0_19_s0), .output_share1(d15_t0_19_s1));
  reg_module u_reg_t0_20_d15 (.clk(clk), .input_share0(d14_t0_20_s0), .input_share1(d14_t0_20_s1), .output_share0(d15_t0_20_s0), .output_share1(d15_t0_20_s1));
  reg_module u_reg_t0_21_d15 (.clk(clk), .input_share0(d14_t0_21_s0), .input_share1(d14_t0_21_s1), .output_share0(d15_t0_21_s0), .output_share1(d15_t0_21_s1));
  reg_module u_reg_t0_22_d15 (.clk(clk), .input_share0(d14_t0_22_s0), .input_share1(d14_t0_22_s1), .output_share0(d15_t0_22_s0), .output_share1(d15_t0_22_s1));
  reg_module u_reg_t0_23_d15 (.clk(clk), .input_share0(d14_t0_23_s0), .input_share1(d14_t0_23_s1), .output_share0(d15_t0_23_s0), .output_share1(d15_t0_23_s1));
  reg_module u_reg_t0_24_d15 (.clk(clk), .input_share0(d14_t0_24_s0), .input_share1(d14_t0_24_s1), .output_share0(d15_t0_24_s0), .output_share1(d15_t0_24_s1));
  reg_module u_reg_t0_25_d15 (.clk(clk), .input_share0(d14_t0_25_s0), .input_share1(d14_t0_25_s1), .output_share0(d15_t0_25_s0), .output_share1(d15_t0_25_s1));
  reg_module u_reg_t0_26_d15 (.clk(clk), .input_share0(d14_t0_26_s0), .input_share1(d14_t0_26_s1), .output_share0(d15_t0_26_s0), .output_share1(d15_t0_26_s1));
  reg_module u_reg_t0_27_d15 (.clk(clk), .input_share0(d14_t0_27_s0), .input_share1(d14_t0_27_s1), .output_share0(d15_t0_27_s0), .output_share1(d15_t0_27_s1));
  reg_module u_reg_t0_28_d15 (.clk(clk), .input_share0(d14_t0_28_s0), .input_share1(d14_t0_28_s1), .output_share0(d15_t0_28_s0), .output_share1(d15_t0_28_s1));
  reg_module u_reg_t0_29_d15 (.clk(clk), .input_share0(d14_t0_29_s0), .input_share1(d14_t0_29_s1), .output_share0(d15_t0_29_s0), .output_share1(d15_t0_29_s1));
  reg_module u_reg_t0_30_d15 (.clk(clk), .input_share0(d14_t0_30_s0), .input_share1(d14_t0_30_s1), .output_share0(d15_t0_30_s0), .output_share1(d15_t0_30_s1));
  reg_module u_reg_t0_31_d15 (.clk(clk), .input_share0(d14_t0_31_s0), .input_share1(d14_t0_31_s1), .output_share0(d15_t0_31_s0), .output_share1(d15_t0_31_s1));
  xor_module u_xor_c15_d15 (.x_share0(d15_i14_s0), .x_share1(d15_i14_s1), .y_share0(d15_t2_14_s0), .y_share1(d15_t2_14_s1), .z_share0(d15_c15_s0), .z_share1(d15_c15_s1));
  xor_module u_xor_o15_d15 (.x_share0(d15_t0_15_s0), .x_share1(d15_t0_15_s1), .y_share0(d15_c15_s0), .y_share1(d15_c15_s1), .z_share0(d15_o15_s0), .z_share1(d15_o15_s1));
  xor_module u_xor_t1_15_d15 (.x_share0(d15_i15_s0), .x_share1(d15_i15_s1), .y_share0(d15_c15_s0), .y_share1(d15_c15_s1), .z_share0(d15_t1_15_s0), .z_share1(d15_t1_15_s1));
  and_module u_and_t2_14_d15 (.clk(clk), .x_share0(d14_t0_14_s0), .x_share1(d14_t0_14_s1), .y_share0(d14_t1_14_s0), .y_share1(d14_t1_14_s1), .rand(r_t2_14), .z_share0(d15_t2_14_s0), .z_share1(d15_t2_14_s1));
  assign r_t2_14 = stage15_share0[0];
  reg_module u_reg_i15_d16 (.clk(clk), .input_share0(d15_i15_s0), .input_share1(d15_i15_s1), .output_share0(d16_i15_s0), .output_share1(d16_i15_s1));
  reg_module u_reg_i16_d16 (.clk(clk), .input_share0(d15_i16_s0), .input_share1(d15_i16_s1), .output_share0(d16_i16_s0), .output_share1(d16_i16_s1));
  reg_module u_reg_i17_d16 (.clk(clk), .input_share0(d15_i17_s0), .input_share1(d15_i17_s1), .output_share0(d16_i17_s0), .output_share1(d16_i17_s1));
  reg_module u_reg_i18_d16 (.clk(clk), .input_share0(d15_i18_s0), .input_share1(d15_i18_s1), .output_share0(d16_i18_s0), .output_share1(d16_i18_s1));
  reg_module u_reg_i19_d16 (.clk(clk), .input_share0(d15_i19_s0), .input_share1(d15_i19_s1), .output_share0(d16_i19_s0), .output_share1(d16_i19_s1));
  reg_module u_reg_i20_d16 (.clk(clk), .input_share0(d15_i20_s0), .input_share1(d15_i20_s1), .output_share0(d16_i20_s0), .output_share1(d16_i20_s1));
  reg_module u_reg_i21_d16 (.clk(clk), .input_share0(d15_i21_s0), .input_share1(d15_i21_s1), .output_share0(d16_i21_s0), .output_share1(d16_i21_s1));
  reg_module u_reg_i22_d16 (.clk(clk), .input_share0(d15_i22_s0), .input_share1(d15_i22_s1), .output_share0(d16_i22_s0), .output_share1(d16_i22_s1));
  reg_module u_reg_i23_d16 (.clk(clk), .input_share0(d15_i23_s0), .input_share1(d15_i23_s1), .output_share0(d16_i23_s0), .output_share1(d16_i23_s1));
  reg_module u_reg_i24_d16 (.clk(clk), .input_share0(d15_i24_s0), .input_share1(d15_i24_s1), .output_share0(d16_i24_s0), .output_share1(d16_i24_s1));
  reg_module u_reg_i25_d16 (.clk(clk), .input_share0(d15_i25_s0), .input_share1(d15_i25_s1), .output_share0(d16_i25_s0), .output_share1(d16_i25_s1));
  reg_module u_reg_i26_d16 (.clk(clk), .input_share0(d15_i26_s0), .input_share1(d15_i26_s1), .output_share0(d16_i26_s0), .output_share1(d16_i26_s1));
  reg_module u_reg_i27_d16 (.clk(clk), .input_share0(d15_i27_s0), .input_share1(d15_i27_s1), .output_share0(d16_i27_s0), .output_share1(d16_i27_s1));
  reg_module u_reg_i28_d16 (.clk(clk), .input_share0(d15_i28_s0), .input_share1(d15_i28_s1), .output_share0(d16_i28_s0), .output_share1(d16_i28_s1));
  reg_module u_reg_i29_d16 (.clk(clk), .input_share0(d15_i29_s0), .input_share1(d15_i29_s1), .output_share0(d16_i29_s0), .output_share1(d16_i29_s1));
  reg_module u_reg_i30_d16 (.clk(clk), .input_share0(d15_i30_s0), .input_share1(d15_i30_s1), .output_share0(d16_i30_s0), .output_share1(d16_i30_s1));
  reg_module u_reg_t0_16_d16 (.clk(clk), .input_share0(d15_t0_16_s0), .input_share1(d15_t0_16_s1), .output_share0(d16_t0_16_s0), .output_share1(d16_t0_16_s1));
  reg_module u_reg_t0_17_d16 (.clk(clk), .input_share0(d15_t0_17_s0), .input_share1(d15_t0_17_s1), .output_share0(d16_t0_17_s0), .output_share1(d16_t0_17_s1));
  reg_module u_reg_t0_18_d16 (.clk(clk), .input_share0(d15_t0_18_s0), .input_share1(d15_t0_18_s1), .output_share0(d16_t0_18_s0), .output_share1(d16_t0_18_s1));
  reg_module u_reg_t0_19_d16 (.clk(clk), .input_share0(d15_t0_19_s0), .input_share1(d15_t0_19_s1), .output_share0(d16_t0_19_s0), .output_share1(d16_t0_19_s1));
  reg_module u_reg_t0_20_d16 (.clk(clk), .input_share0(d15_t0_20_s0), .input_share1(d15_t0_20_s1), .output_share0(d16_t0_20_s0), .output_share1(d16_t0_20_s1));
  reg_module u_reg_t0_21_d16 (.clk(clk), .input_share0(d15_t0_21_s0), .input_share1(d15_t0_21_s1), .output_share0(d16_t0_21_s0), .output_share1(d16_t0_21_s1));
  reg_module u_reg_t0_22_d16 (.clk(clk), .input_share0(d15_t0_22_s0), .input_share1(d15_t0_22_s1), .output_share0(d16_t0_22_s0), .output_share1(d16_t0_22_s1));
  reg_module u_reg_t0_23_d16 (.clk(clk), .input_share0(d15_t0_23_s0), .input_share1(d15_t0_23_s1), .output_share0(d16_t0_23_s0), .output_share1(d16_t0_23_s1));
  reg_module u_reg_t0_24_d16 (.clk(clk), .input_share0(d15_t0_24_s0), .input_share1(d15_t0_24_s1), .output_share0(d16_t0_24_s0), .output_share1(d16_t0_24_s1));
  reg_module u_reg_t0_25_d16 (.clk(clk), .input_share0(d15_t0_25_s0), .input_share1(d15_t0_25_s1), .output_share0(d16_t0_25_s0), .output_share1(d16_t0_25_s1));
  reg_module u_reg_t0_26_d16 (.clk(clk), .input_share0(d15_t0_26_s0), .input_share1(d15_t0_26_s1), .output_share0(d16_t0_26_s0), .output_share1(d16_t0_26_s1));
  reg_module u_reg_t0_27_d16 (.clk(clk), .input_share0(d15_t0_27_s0), .input_share1(d15_t0_27_s1), .output_share0(d16_t0_27_s0), .output_share1(d16_t0_27_s1));
  reg_module u_reg_t0_28_d16 (.clk(clk), .input_share0(d15_t0_28_s0), .input_share1(d15_t0_28_s1), .output_share0(d16_t0_28_s0), .output_share1(d16_t0_28_s1));
  reg_module u_reg_t0_29_d16 (.clk(clk), .input_share0(d15_t0_29_s0), .input_share1(d15_t0_29_s1), .output_share0(d16_t0_29_s0), .output_share1(d16_t0_29_s1));
  reg_module u_reg_t0_30_d16 (.clk(clk), .input_share0(d15_t0_30_s0), .input_share1(d15_t0_30_s1), .output_share0(d16_t0_30_s0), .output_share1(d16_t0_30_s1));
  reg_module u_reg_t0_31_d16 (.clk(clk), .input_share0(d15_t0_31_s0), .input_share1(d15_t0_31_s1), .output_share0(d16_t0_31_s0), .output_share1(d16_t0_31_s1));
  xor_module u_xor_c16_d16 (.x_share0(d16_i15_s0), .x_share1(d16_i15_s1), .y_share0(d16_t2_15_s0), .y_share1(d16_t2_15_s1), .z_share0(d16_c16_s0), .z_share1(d16_c16_s1));
  xor_module u_xor_o16_d16 (.x_share0(d16_t0_16_s0), .x_share1(d16_t0_16_s1), .y_share0(d16_c16_s0), .y_share1(d16_c16_s1), .z_share0(d16_o16_s0), .z_share1(d16_o16_s1));
  xor_module u_xor_t1_16_d16 (.x_share0(d16_i16_s0), .x_share1(d16_i16_s1), .y_share0(d16_c16_s0), .y_share1(d16_c16_s1), .z_share0(d16_t1_16_s0), .z_share1(d16_t1_16_s1));
  and_module u_and_t2_15_d16 (.clk(clk), .x_share0(d15_t0_15_s0), .x_share1(d15_t0_15_s1), .y_share0(d15_t1_15_s0), .y_share1(d15_t1_15_s1), .rand(r_t2_15), .z_share0(d16_t2_15_s0), .z_share1(d16_t2_15_s1));
  assign r_t2_15 = stage16_share0[1];
  reg_module u_reg_i16_d17 (.clk(clk), .input_share0(d16_i16_s0), .input_share1(d16_i16_s1), .output_share0(d17_i16_s0), .output_share1(d17_i16_s1));
  reg_module u_reg_i17_d17 (.clk(clk), .input_share0(d16_i17_s0), .input_share1(d16_i17_s1), .output_share0(d17_i17_s0), .output_share1(d17_i17_s1));
  reg_module u_reg_i18_d17 (.clk(clk), .input_share0(d16_i18_s0), .input_share1(d16_i18_s1), .output_share0(d17_i18_s0), .output_share1(d17_i18_s1));
  reg_module u_reg_i19_d17 (.clk(clk), .input_share0(d16_i19_s0), .input_share1(d16_i19_s1), .output_share0(d17_i19_s0), .output_share1(d17_i19_s1));
  reg_module u_reg_i20_d17 (.clk(clk), .input_share0(d16_i20_s0), .input_share1(d16_i20_s1), .output_share0(d17_i20_s0), .output_share1(d17_i20_s1));
  reg_module u_reg_i21_d17 (.clk(clk), .input_share0(d16_i21_s0), .input_share1(d16_i21_s1), .output_share0(d17_i21_s0), .output_share1(d17_i21_s1));
  reg_module u_reg_i22_d17 (.clk(clk), .input_share0(d16_i22_s0), .input_share1(d16_i22_s1), .output_share0(d17_i22_s0), .output_share1(d17_i22_s1));
  reg_module u_reg_i23_d17 (.clk(clk), .input_share0(d16_i23_s0), .input_share1(d16_i23_s1), .output_share0(d17_i23_s0), .output_share1(d17_i23_s1));
  reg_module u_reg_i24_d17 (.clk(clk), .input_share0(d16_i24_s0), .input_share1(d16_i24_s1), .output_share0(d17_i24_s0), .output_share1(d17_i24_s1));
  reg_module u_reg_i25_d17 (.clk(clk), .input_share0(d16_i25_s0), .input_share1(d16_i25_s1), .output_share0(d17_i25_s0), .output_share1(d17_i25_s1));
  reg_module u_reg_i26_d17 (.clk(clk), .input_share0(d16_i26_s0), .input_share1(d16_i26_s1), .output_share0(d17_i26_s0), .output_share1(d17_i26_s1));
  reg_module u_reg_i27_d17 (.clk(clk), .input_share0(d16_i27_s0), .input_share1(d16_i27_s1), .output_share0(d17_i27_s0), .output_share1(d17_i27_s1));
  reg_module u_reg_i28_d17 (.clk(clk), .input_share0(d16_i28_s0), .input_share1(d16_i28_s1), .output_share0(d17_i28_s0), .output_share1(d17_i28_s1));
  reg_module u_reg_i29_d17 (.clk(clk), .input_share0(d16_i29_s0), .input_share1(d16_i29_s1), .output_share0(d17_i29_s0), .output_share1(d17_i29_s1));
  reg_module u_reg_i30_d17 (.clk(clk), .input_share0(d16_i30_s0), .input_share1(d16_i30_s1), .output_share0(d17_i30_s0), .output_share1(d17_i30_s1));
  reg_module u_reg_t0_17_d17 (.clk(clk), .input_share0(d16_t0_17_s0), .input_share1(d16_t0_17_s1), .output_share0(d17_t0_17_s0), .output_share1(d17_t0_17_s1));
  reg_module u_reg_t0_18_d17 (.clk(clk), .input_share0(d16_t0_18_s0), .input_share1(d16_t0_18_s1), .output_share0(d17_t0_18_s0), .output_share1(d17_t0_18_s1));
  reg_module u_reg_t0_19_d17 (.clk(clk), .input_share0(d16_t0_19_s0), .input_share1(d16_t0_19_s1), .output_share0(d17_t0_19_s0), .output_share1(d17_t0_19_s1));
  reg_module u_reg_t0_20_d17 (.clk(clk), .input_share0(d16_t0_20_s0), .input_share1(d16_t0_20_s1), .output_share0(d17_t0_20_s0), .output_share1(d17_t0_20_s1));
  reg_module u_reg_t0_21_d17 (.clk(clk), .input_share0(d16_t0_21_s0), .input_share1(d16_t0_21_s1), .output_share0(d17_t0_21_s0), .output_share1(d17_t0_21_s1));
  reg_module u_reg_t0_22_d17 (.clk(clk), .input_share0(d16_t0_22_s0), .input_share1(d16_t0_22_s1), .output_share0(d17_t0_22_s0), .output_share1(d17_t0_22_s1));
  reg_module u_reg_t0_23_d17 (.clk(clk), .input_share0(d16_t0_23_s0), .input_share1(d16_t0_23_s1), .output_share0(d17_t0_23_s0), .output_share1(d17_t0_23_s1));
  reg_module u_reg_t0_24_d17 (.clk(clk), .input_share0(d16_t0_24_s0), .input_share1(d16_t0_24_s1), .output_share0(d17_t0_24_s0), .output_share1(d17_t0_24_s1));
  reg_module u_reg_t0_25_d17 (.clk(clk), .input_share0(d16_t0_25_s0), .input_share1(d16_t0_25_s1), .output_share0(d17_t0_25_s0), .output_share1(d17_t0_25_s1));
  reg_module u_reg_t0_26_d17 (.clk(clk), .input_share0(d16_t0_26_s0), .input_share1(d16_t0_26_s1), .output_share0(d17_t0_26_s0), .output_share1(d17_t0_26_s1));
  reg_module u_reg_t0_27_d17 (.clk(clk), .input_share0(d16_t0_27_s0), .input_share1(d16_t0_27_s1), .output_share0(d17_t0_27_s0), .output_share1(d17_t0_27_s1));
  reg_module u_reg_t0_28_d17 (.clk(clk), .input_share0(d16_t0_28_s0), .input_share1(d16_t0_28_s1), .output_share0(d17_t0_28_s0), .output_share1(d17_t0_28_s1));
  reg_module u_reg_t0_29_d17 (.clk(clk), .input_share0(d16_t0_29_s0), .input_share1(d16_t0_29_s1), .output_share0(d17_t0_29_s0), .output_share1(d17_t0_29_s1));
  reg_module u_reg_t0_30_d17 (.clk(clk), .input_share0(d16_t0_30_s0), .input_share1(d16_t0_30_s1), .output_share0(d17_t0_30_s0), .output_share1(d17_t0_30_s1));
  reg_module u_reg_t0_31_d17 (.clk(clk), .input_share0(d16_t0_31_s0), .input_share1(d16_t0_31_s1), .output_share0(d17_t0_31_s0), .output_share1(d17_t0_31_s1));
  xor_module u_xor_c17_d17 (.x_share0(d17_i16_s0), .x_share1(d17_i16_s1), .y_share0(d17_t2_16_s0), .y_share1(d17_t2_16_s1), .z_share0(d17_c17_s0), .z_share1(d17_c17_s1));
  xor_module u_xor_o17_d17 (.x_share0(d17_t0_17_s0), .x_share1(d17_t0_17_s1), .y_share0(d17_c17_s0), .y_share1(d17_c17_s1), .z_share0(d17_o17_s0), .z_share1(d17_o17_s1));
  xor_module u_xor_t1_17_d17 (.x_share0(d17_i17_s0), .x_share1(d17_i17_s1), .y_share0(d17_c17_s0), .y_share1(d17_c17_s1), .z_share0(d17_t1_17_s0), .z_share1(d17_t1_17_s1));
  and_module u_and_t2_16_d17 (.clk(clk), .x_share0(d16_t0_16_s0), .x_share1(d16_t0_16_s1), .y_share0(d16_t1_16_s0), .y_share1(d16_t1_16_s1), .rand(r_t2_16), .z_share0(d17_t2_16_s0), .z_share1(d17_t2_16_s1));
  assign r_t2_16 = stage17_share0[2];
  reg_module u_reg_i17_d18 (.clk(clk), .input_share0(d17_i17_s0), .input_share1(d17_i17_s1), .output_share0(d18_i17_s0), .output_share1(d18_i17_s1));
  reg_module u_reg_i18_d18 (.clk(clk), .input_share0(d17_i18_s0), .input_share1(d17_i18_s1), .output_share0(d18_i18_s0), .output_share1(d18_i18_s1));
  reg_module u_reg_i19_d18 (.clk(clk), .input_share0(d17_i19_s0), .input_share1(d17_i19_s1), .output_share0(d18_i19_s0), .output_share1(d18_i19_s1));
  reg_module u_reg_i20_d18 (.clk(clk), .input_share0(d17_i20_s0), .input_share1(d17_i20_s1), .output_share0(d18_i20_s0), .output_share1(d18_i20_s1));
  reg_module u_reg_i21_d18 (.clk(clk), .input_share0(d17_i21_s0), .input_share1(d17_i21_s1), .output_share0(d18_i21_s0), .output_share1(d18_i21_s1));
  reg_module u_reg_i22_d18 (.clk(clk), .input_share0(d17_i22_s0), .input_share1(d17_i22_s1), .output_share0(d18_i22_s0), .output_share1(d18_i22_s1));
  reg_module u_reg_i23_d18 (.clk(clk), .input_share0(d17_i23_s0), .input_share1(d17_i23_s1), .output_share0(d18_i23_s0), .output_share1(d18_i23_s1));
  reg_module u_reg_i24_d18 (.clk(clk), .input_share0(d17_i24_s0), .input_share1(d17_i24_s1), .output_share0(d18_i24_s0), .output_share1(d18_i24_s1));
  reg_module u_reg_i25_d18 (.clk(clk), .input_share0(d17_i25_s0), .input_share1(d17_i25_s1), .output_share0(d18_i25_s0), .output_share1(d18_i25_s1));
  reg_module u_reg_i26_d18 (.clk(clk), .input_share0(d17_i26_s0), .input_share1(d17_i26_s1), .output_share0(d18_i26_s0), .output_share1(d18_i26_s1));
  reg_module u_reg_i27_d18 (.clk(clk), .input_share0(d17_i27_s0), .input_share1(d17_i27_s1), .output_share0(d18_i27_s0), .output_share1(d18_i27_s1));
  reg_module u_reg_i28_d18 (.clk(clk), .input_share0(d17_i28_s0), .input_share1(d17_i28_s1), .output_share0(d18_i28_s0), .output_share1(d18_i28_s1));
  reg_module u_reg_i29_d18 (.clk(clk), .input_share0(d17_i29_s0), .input_share1(d17_i29_s1), .output_share0(d18_i29_s0), .output_share1(d18_i29_s1));
  reg_module u_reg_i30_d18 (.clk(clk), .input_share0(d17_i30_s0), .input_share1(d17_i30_s1), .output_share0(d18_i30_s0), .output_share1(d18_i30_s1));
  reg_module u_reg_t0_18_d18 (.clk(clk), .input_share0(d17_t0_18_s0), .input_share1(d17_t0_18_s1), .output_share0(d18_t0_18_s0), .output_share1(d18_t0_18_s1));
  reg_module u_reg_t0_19_d18 (.clk(clk), .input_share0(d17_t0_19_s0), .input_share1(d17_t0_19_s1), .output_share0(d18_t0_19_s0), .output_share1(d18_t0_19_s1));
  reg_module u_reg_t0_20_d18 (.clk(clk), .input_share0(d17_t0_20_s0), .input_share1(d17_t0_20_s1), .output_share0(d18_t0_20_s0), .output_share1(d18_t0_20_s1));
  reg_module u_reg_t0_21_d18 (.clk(clk), .input_share0(d17_t0_21_s0), .input_share1(d17_t0_21_s1), .output_share0(d18_t0_21_s0), .output_share1(d18_t0_21_s1));
  reg_module u_reg_t0_22_d18 (.clk(clk), .input_share0(d17_t0_22_s0), .input_share1(d17_t0_22_s1), .output_share0(d18_t0_22_s0), .output_share1(d18_t0_22_s1));
  reg_module u_reg_t0_23_d18 (.clk(clk), .input_share0(d17_t0_23_s0), .input_share1(d17_t0_23_s1), .output_share0(d18_t0_23_s0), .output_share1(d18_t0_23_s1));
  reg_module u_reg_t0_24_d18 (.clk(clk), .input_share0(d17_t0_24_s0), .input_share1(d17_t0_24_s1), .output_share0(d18_t0_24_s0), .output_share1(d18_t0_24_s1));
  reg_module u_reg_t0_25_d18 (.clk(clk), .input_share0(d17_t0_25_s0), .input_share1(d17_t0_25_s1), .output_share0(d18_t0_25_s0), .output_share1(d18_t0_25_s1));
  reg_module u_reg_t0_26_d18 (.clk(clk), .input_share0(d17_t0_26_s0), .input_share1(d17_t0_26_s1), .output_share0(d18_t0_26_s0), .output_share1(d18_t0_26_s1));
  reg_module u_reg_t0_27_d18 (.clk(clk), .input_share0(d17_t0_27_s0), .input_share1(d17_t0_27_s1), .output_share0(d18_t0_27_s0), .output_share1(d18_t0_27_s1));
  reg_module u_reg_t0_28_d18 (.clk(clk), .input_share0(d17_t0_28_s0), .input_share1(d17_t0_28_s1), .output_share0(d18_t0_28_s0), .output_share1(d18_t0_28_s1));
  reg_module u_reg_t0_29_d18 (.clk(clk), .input_share0(d17_t0_29_s0), .input_share1(d17_t0_29_s1), .output_share0(d18_t0_29_s0), .output_share1(d18_t0_29_s1));
  reg_module u_reg_t0_30_d18 (.clk(clk), .input_share0(d17_t0_30_s0), .input_share1(d17_t0_30_s1), .output_share0(d18_t0_30_s0), .output_share1(d18_t0_30_s1));
  reg_module u_reg_t0_31_d18 (.clk(clk), .input_share0(d17_t0_31_s0), .input_share1(d17_t0_31_s1), .output_share0(d18_t0_31_s0), .output_share1(d18_t0_31_s1));
  xor_module u_xor_c18_d18 (.x_share0(d18_i17_s0), .x_share1(d18_i17_s1), .y_share0(d18_t2_17_s0), .y_share1(d18_t2_17_s1), .z_share0(d18_c18_s0), .z_share1(d18_c18_s1));
  xor_module u_xor_o18_d18 (.x_share0(d18_t0_18_s0), .x_share1(d18_t0_18_s1), .y_share0(d18_c18_s0), .y_share1(d18_c18_s1), .z_share0(d18_o18_s0), .z_share1(d18_o18_s1));
  xor_module u_xor_t1_18_d18 (.x_share0(d18_i18_s0), .x_share1(d18_i18_s1), .y_share0(d18_c18_s0), .y_share1(d18_c18_s1), .z_share0(d18_t1_18_s0), .z_share1(d18_t1_18_s1));
  and_module u_and_t2_17_d18 (.clk(clk), .x_share0(d17_t0_17_s0), .x_share1(d17_t0_17_s1), .y_share0(d17_t1_17_s0), .y_share1(d17_t1_17_s1), .rand(r_t2_17), .z_share0(d18_t2_17_s0), .z_share1(d18_t2_17_s1));
  assign r_t2_17 = stage18_share0[0];
  reg_module u_reg_i18_d19 (.clk(clk), .input_share0(d18_i18_s0), .input_share1(d18_i18_s1), .output_share0(d19_i18_s0), .output_share1(d19_i18_s1));
  reg_module u_reg_i19_d19 (.clk(clk), .input_share0(d18_i19_s0), .input_share1(d18_i19_s1), .output_share0(d19_i19_s0), .output_share1(d19_i19_s1));
  reg_module u_reg_i20_d19 (.clk(clk), .input_share0(d18_i20_s0), .input_share1(d18_i20_s1), .output_share0(d19_i20_s0), .output_share1(d19_i20_s1));
  reg_module u_reg_i21_d19 (.clk(clk), .input_share0(d18_i21_s0), .input_share1(d18_i21_s1), .output_share0(d19_i21_s0), .output_share1(d19_i21_s1));
  reg_module u_reg_i22_d19 (.clk(clk), .input_share0(d18_i22_s0), .input_share1(d18_i22_s1), .output_share0(d19_i22_s0), .output_share1(d19_i22_s1));
  reg_module u_reg_i23_d19 (.clk(clk), .input_share0(d18_i23_s0), .input_share1(d18_i23_s1), .output_share0(d19_i23_s0), .output_share1(d19_i23_s1));
  reg_module u_reg_i24_d19 (.clk(clk), .input_share0(d18_i24_s0), .input_share1(d18_i24_s1), .output_share0(d19_i24_s0), .output_share1(d19_i24_s1));
  reg_module u_reg_i25_d19 (.clk(clk), .input_share0(d18_i25_s0), .input_share1(d18_i25_s1), .output_share0(d19_i25_s0), .output_share1(d19_i25_s1));
  reg_module u_reg_i26_d19 (.clk(clk), .input_share0(d18_i26_s0), .input_share1(d18_i26_s1), .output_share0(d19_i26_s0), .output_share1(d19_i26_s1));
  reg_module u_reg_i27_d19 (.clk(clk), .input_share0(d18_i27_s0), .input_share1(d18_i27_s1), .output_share0(d19_i27_s0), .output_share1(d19_i27_s1));
  reg_module u_reg_i28_d19 (.clk(clk), .input_share0(d18_i28_s0), .input_share1(d18_i28_s1), .output_share0(d19_i28_s0), .output_share1(d19_i28_s1));
  reg_module u_reg_i29_d19 (.clk(clk), .input_share0(d18_i29_s0), .input_share1(d18_i29_s1), .output_share0(d19_i29_s0), .output_share1(d19_i29_s1));
  reg_module u_reg_i30_d19 (.clk(clk), .input_share0(d18_i30_s0), .input_share1(d18_i30_s1), .output_share0(d19_i30_s0), .output_share1(d19_i30_s1));
  reg_module u_reg_t0_19_d19 (.clk(clk), .input_share0(d18_t0_19_s0), .input_share1(d18_t0_19_s1), .output_share0(d19_t0_19_s0), .output_share1(d19_t0_19_s1));
  reg_module u_reg_t0_20_d19 (.clk(clk), .input_share0(d18_t0_20_s0), .input_share1(d18_t0_20_s1), .output_share0(d19_t0_20_s0), .output_share1(d19_t0_20_s1));
  reg_module u_reg_t0_21_d19 (.clk(clk), .input_share0(d18_t0_21_s0), .input_share1(d18_t0_21_s1), .output_share0(d19_t0_21_s0), .output_share1(d19_t0_21_s1));
  reg_module u_reg_t0_22_d19 (.clk(clk), .input_share0(d18_t0_22_s0), .input_share1(d18_t0_22_s1), .output_share0(d19_t0_22_s0), .output_share1(d19_t0_22_s1));
  reg_module u_reg_t0_23_d19 (.clk(clk), .input_share0(d18_t0_23_s0), .input_share1(d18_t0_23_s1), .output_share0(d19_t0_23_s0), .output_share1(d19_t0_23_s1));
  reg_module u_reg_t0_24_d19 (.clk(clk), .input_share0(d18_t0_24_s0), .input_share1(d18_t0_24_s1), .output_share0(d19_t0_24_s0), .output_share1(d19_t0_24_s1));
  reg_module u_reg_t0_25_d19 (.clk(clk), .input_share0(d18_t0_25_s0), .input_share1(d18_t0_25_s1), .output_share0(d19_t0_25_s0), .output_share1(d19_t0_25_s1));
  reg_module u_reg_t0_26_d19 (.clk(clk), .input_share0(d18_t0_26_s0), .input_share1(d18_t0_26_s1), .output_share0(d19_t0_26_s0), .output_share1(d19_t0_26_s1));
  reg_module u_reg_t0_27_d19 (.clk(clk), .input_share0(d18_t0_27_s0), .input_share1(d18_t0_27_s1), .output_share0(d19_t0_27_s0), .output_share1(d19_t0_27_s1));
  reg_module u_reg_t0_28_d19 (.clk(clk), .input_share0(d18_t0_28_s0), .input_share1(d18_t0_28_s1), .output_share0(d19_t0_28_s0), .output_share1(d19_t0_28_s1));
  reg_module u_reg_t0_29_d19 (.clk(clk), .input_share0(d18_t0_29_s0), .input_share1(d18_t0_29_s1), .output_share0(d19_t0_29_s0), .output_share1(d19_t0_29_s1));
  reg_module u_reg_t0_30_d19 (.clk(clk), .input_share0(d18_t0_30_s0), .input_share1(d18_t0_30_s1), .output_share0(d19_t0_30_s0), .output_share1(d19_t0_30_s1));
  reg_module u_reg_t0_31_d19 (.clk(clk), .input_share0(d18_t0_31_s0), .input_share1(d18_t0_31_s1), .output_share0(d19_t0_31_s0), .output_share1(d19_t0_31_s1));
  xor_module u_xor_c19_d19 (.x_share0(d19_i18_s0), .x_share1(d19_i18_s1), .y_share0(d19_t2_18_s0), .y_share1(d19_t2_18_s1), .z_share0(d19_c19_s0), .z_share1(d19_c19_s1));
  xor_module u_xor_o19_d19 (.x_share0(d19_t0_19_s0), .x_share1(d19_t0_19_s1), .y_share0(d19_c19_s0), .y_share1(d19_c19_s1), .z_share0(d19_o19_s0), .z_share1(d19_o19_s1));
  xor_module u_xor_t1_19_d19 (.x_share0(d19_i19_s0), .x_share1(d19_i19_s1), .y_share0(d19_c19_s0), .y_share1(d19_c19_s1), .z_share0(d19_t1_19_s0), .z_share1(d19_t1_19_s1));
  and_module u_and_t2_18_d19 (.clk(clk), .x_share0(d18_t0_18_s0), .x_share1(d18_t0_18_s1), .y_share0(d18_t1_18_s0), .y_share1(d18_t1_18_s1), .rand(r_t2_18), .z_share0(d19_t2_18_s0), .z_share1(d19_t2_18_s1));
  assign r_t2_18 = stage19_share0[1];
  reg_module u_reg_i19_d20 (.clk(clk), .input_share0(d19_i19_s0), .input_share1(d19_i19_s1), .output_share0(d20_i19_s0), .output_share1(d20_i19_s1));
  reg_module u_reg_i20_d20 (.clk(clk), .input_share0(d19_i20_s0), .input_share1(d19_i20_s1), .output_share0(d20_i20_s0), .output_share1(d20_i20_s1));
  reg_module u_reg_i21_d20 (.clk(clk), .input_share0(d19_i21_s0), .input_share1(d19_i21_s1), .output_share0(d20_i21_s0), .output_share1(d20_i21_s1));
  reg_module u_reg_i22_d20 (.clk(clk), .input_share0(d19_i22_s0), .input_share1(d19_i22_s1), .output_share0(d20_i22_s0), .output_share1(d20_i22_s1));
  reg_module u_reg_i23_d20 (.clk(clk), .input_share0(d19_i23_s0), .input_share1(d19_i23_s1), .output_share0(d20_i23_s0), .output_share1(d20_i23_s1));
  reg_module u_reg_i24_d20 (.clk(clk), .input_share0(d19_i24_s0), .input_share1(d19_i24_s1), .output_share0(d20_i24_s0), .output_share1(d20_i24_s1));
  reg_module u_reg_i25_d20 (.clk(clk), .input_share0(d19_i25_s0), .input_share1(d19_i25_s1), .output_share0(d20_i25_s0), .output_share1(d20_i25_s1));
  reg_module u_reg_i26_d20 (.clk(clk), .input_share0(d19_i26_s0), .input_share1(d19_i26_s1), .output_share0(d20_i26_s0), .output_share1(d20_i26_s1));
  reg_module u_reg_i27_d20 (.clk(clk), .input_share0(d19_i27_s0), .input_share1(d19_i27_s1), .output_share0(d20_i27_s0), .output_share1(d20_i27_s1));
  reg_module u_reg_i28_d20 (.clk(clk), .input_share0(d19_i28_s0), .input_share1(d19_i28_s1), .output_share0(d20_i28_s0), .output_share1(d20_i28_s1));
  reg_module u_reg_i29_d20 (.clk(clk), .input_share0(d19_i29_s0), .input_share1(d19_i29_s1), .output_share0(d20_i29_s0), .output_share1(d20_i29_s1));
  reg_module u_reg_i30_d20 (.clk(clk), .input_share0(d19_i30_s0), .input_share1(d19_i30_s1), .output_share0(d20_i30_s0), .output_share1(d20_i30_s1));
  reg_module u_reg_t0_20_d20 (.clk(clk), .input_share0(d19_t0_20_s0), .input_share1(d19_t0_20_s1), .output_share0(d20_t0_20_s0), .output_share1(d20_t0_20_s1));
  reg_module u_reg_t0_21_d20 (.clk(clk), .input_share0(d19_t0_21_s0), .input_share1(d19_t0_21_s1), .output_share0(d20_t0_21_s0), .output_share1(d20_t0_21_s1));
  reg_module u_reg_t0_22_d20 (.clk(clk), .input_share0(d19_t0_22_s0), .input_share1(d19_t0_22_s1), .output_share0(d20_t0_22_s0), .output_share1(d20_t0_22_s1));
  reg_module u_reg_t0_23_d20 (.clk(clk), .input_share0(d19_t0_23_s0), .input_share1(d19_t0_23_s1), .output_share0(d20_t0_23_s0), .output_share1(d20_t0_23_s1));
  reg_module u_reg_t0_24_d20 (.clk(clk), .input_share0(d19_t0_24_s0), .input_share1(d19_t0_24_s1), .output_share0(d20_t0_24_s0), .output_share1(d20_t0_24_s1));
  reg_module u_reg_t0_25_d20 (.clk(clk), .input_share0(d19_t0_25_s0), .input_share1(d19_t0_25_s1), .output_share0(d20_t0_25_s0), .output_share1(d20_t0_25_s1));
  reg_module u_reg_t0_26_d20 (.clk(clk), .input_share0(d19_t0_26_s0), .input_share1(d19_t0_26_s1), .output_share0(d20_t0_26_s0), .output_share1(d20_t0_26_s1));
  reg_module u_reg_t0_27_d20 (.clk(clk), .input_share0(d19_t0_27_s0), .input_share1(d19_t0_27_s1), .output_share0(d20_t0_27_s0), .output_share1(d20_t0_27_s1));
  reg_module u_reg_t0_28_d20 (.clk(clk), .input_share0(d19_t0_28_s0), .input_share1(d19_t0_28_s1), .output_share0(d20_t0_28_s0), .output_share1(d20_t0_28_s1));
  reg_module u_reg_t0_29_d20 (.clk(clk), .input_share0(d19_t0_29_s0), .input_share1(d19_t0_29_s1), .output_share0(d20_t0_29_s0), .output_share1(d20_t0_29_s1));
  reg_module u_reg_t0_30_d20 (.clk(clk), .input_share0(d19_t0_30_s0), .input_share1(d19_t0_30_s1), .output_share0(d20_t0_30_s0), .output_share1(d20_t0_30_s1));
  reg_module u_reg_t0_31_d20 (.clk(clk), .input_share0(d19_t0_31_s0), .input_share1(d19_t0_31_s1), .output_share0(d20_t0_31_s0), .output_share1(d20_t0_31_s1));
  xor_module u_xor_c20_d20 (.x_share0(d20_i19_s0), .x_share1(d20_i19_s1), .y_share0(d20_t2_19_s0), .y_share1(d20_t2_19_s1), .z_share0(d20_c20_s0), .z_share1(d20_c20_s1));
  xor_module u_xor_o20_d20 (.x_share0(d20_t0_20_s0), .x_share1(d20_t0_20_s1), .y_share0(d20_c20_s0), .y_share1(d20_c20_s1), .z_share0(d20_o20_s0), .z_share1(d20_o20_s1));
  xor_module u_xor_t1_20_d20 (.x_share0(d20_i20_s0), .x_share1(d20_i20_s1), .y_share0(d20_c20_s0), .y_share1(d20_c20_s1), .z_share0(d20_t1_20_s0), .z_share1(d20_t1_20_s1));
  and_module u_and_t2_19_d20 (.clk(clk), .x_share0(d19_t0_19_s0), .x_share1(d19_t0_19_s1), .y_share0(d19_t1_19_s0), .y_share1(d19_t1_19_s1), .rand(r_t2_19), .z_share0(d20_t2_19_s0), .z_share1(d20_t2_19_s1));
  assign r_t2_19 = stage20_share0[2];
  reg_module u_reg_i20_d21 (.clk(clk), .input_share0(d20_i20_s0), .input_share1(d20_i20_s1), .output_share0(d21_i20_s0), .output_share1(d21_i20_s1));
  reg_module u_reg_i21_d21 (.clk(clk), .input_share0(d20_i21_s0), .input_share1(d20_i21_s1), .output_share0(d21_i21_s0), .output_share1(d21_i21_s1));
  reg_module u_reg_i22_d21 (.clk(clk), .input_share0(d20_i22_s0), .input_share1(d20_i22_s1), .output_share0(d21_i22_s0), .output_share1(d21_i22_s1));
  reg_module u_reg_i23_d21 (.clk(clk), .input_share0(d20_i23_s0), .input_share1(d20_i23_s1), .output_share0(d21_i23_s0), .output_share1(d21_i23_s1));
  reg_module u_reg_i24_d21 (.clk(clk), .input_share0(d20_i24_s0), .input_share1(d20_i24_s1), .output_share0(d21_i24_s0), .output_share1(d21_i24_s1));
  reg_module u_reg_i25_d21 (.clk(clk), .input_share0(d20_i25_s0), .input_share1(d20_i25_s1), .output_share0(d21_i25_s0), .output_share1(d21_i25_s1));
  reg_module u_reg_i26_d21 (.clk(clk), .input_share0(d20_i26_s0), .input_share1(d20_i26_s1), .output_share0(d21_i26_s0), .output_share1(d21_i26_s1));
  reg_module u_reg_i27_d21 (.clk(clk), .input_share0(d20_i27_s0), .input_share1(d20_i27_s1), .output_share0(d21_i27_s0), .output_share1(d21_i27_s1));
  reg_module u_reg_i28_d21 (.clk(clk), .input_share0(d20_i28_s0), .input_share1(d20_i28_s1), .output_share0(d21_i28_s0), .output_share1(d21_i28_s1));
  reg_module u_reg_i29_d21 (.clk(clk), .input_share0(d20_i29_s0), .input_share1(d20_i29_s1), .output_share0(d21_i29_s0), .output_share1(d21_i29_s1));
  reg_module u_reg_i30_d21 (.clk(clk), .input_share0(d20_i30_s0), .input_share1(d20_i30_s1), .output_share0(d21_i30_s0), .output_share1(d21_i30_s1));
  reg_module u_reg_t0_21_d21 (.clk(clk), .input_share0(d20_t0_21_s0), .input_share1(d20_t0_21_s1), .output_share0(d21_t0_21_s0), .output_share1(d21_t0_21_s1));
  reg_module u_reg_t0_22_d21 (.clk(clk), .input_share0(d20_t0_22_s0), .input_share1(d20_t0_22_s1), .output_share0(d21_t0_22_s0), .output_share1(d21_t0_22_s1));
  reg_module u_reg_t0_23_d21 (.clk(clk), .input_share0(d20_t0_23_s0), .input_share1(d20_t0_23_s1), .output_share0(d21_t0_23_s0), .output_share1(d21_t0_23_s1));
  reg_module u_reg_t0_24_d21 (.clk(clk), .input_share0(d20_t0_24_s0), .input_share1(d20_t0_24_s1), .output_share0(d21_t0_24_s0), .output_share1(d21_t0_24_s1));
  reg_module u_reg_t0_25_d21 (.clk(clk), .input_share0(d20_t0_25_s0), .input_share1(d20_t0_25_s1), .output_share0(d21_t0_25_s0), .output_share1(d21_t0_25_s1));
  reg_module u_reg_t0_26_d21 (.clk(clk), .input_share0(d20_t0_26_s0), .input_share1(d20_t0_26_s1), .output_share0(d21_t0_26_s0), .output_share1(d21_t0_26_s1));
  reg_module u_reg_t0_27_d21 (.clk(clk), .input_share0(d20_t0_27_s0), .input_share1(d20_t0_27_s1), .output_share0(d21_t0_27_s0), .output_share1(d21_t0_27_s1));
  reg_module u_reg_t0_28_d21 (.clk(clk), .input_share0(d20_t0_28_s0), .input_share1(d20_t0_28_s1), .output_share0(d21_t0_28_s0), .output_share1(d21_t0_28_s1));
  reg_module u_reg_t0_29_d21 (.clk(clk), .input_share0(d20_t0_29_s0), .input_share1(d20_t0_29_s1), .output_share0(d21_t0_29_s0), .output_share1(d21_t0_29_s1));
  reg_module u_reg_t0_30_d21 (.clk(clk), .input_share0(d20_t0_30_s0), .input_share1(d20_t0_30_s1), .output_share0(d21_t0_30_s0), .output_share1(d21_t0_30_s1));
  reg_module u_reg_t0_31_d21 (.clk(clk), .input_share0(d20_t0_31_s0), .input_share1(d20_t0_31_s1), .output_share0(d21_t0_31_s0), .output_share1(d21_t0_31_s1));
  xor_module u_xor_c21_d21 (.x_share0(d21_i20_s0), .x_share1(d21_i20_s1), .y_share0(d21_t2_20_s0), .y_share1(d21_t2_20_s1), .z_share0(d21_c21_s0), .z_share1(d21_c21_s1));
  xor_module u_xor_o21_d21 (.x_share0(d21_t0_21_s0), .x_share1(d21_t0_21_s1), .y_share0(d21_c21_s0), .y_share1(d21_c21_s1), .z_share0(d21_o21_s0), .z_share1(d21_o21_s1));
  xor_module u_xor_t1_21_d21 (.x_share0(d21_i21_s0), .x_share1(d21_i21_s1), .y_share0(d21_c21_s0), .y_share1(d21_c21_s1), .z_share0(d21_t1_21_s0), .z_share1(d21_t1_21_s1));
  and_module u_and_t2_20_d21 (.clk(clk), .x_share0(d20_t0_20_s0), .x_share1(d20_t0_20_s1), .y_share0(d20_t1_20_s0), .y_share1(d20_t1_20_s1), .rand(r_t2_20), .z_share0(d21_t2_20_s0), .z_share1(d21_t2_20_s1));
  assign r_t2_20 = stage21_share0[0];
  reg_module u_reg_i21_d22 (.clk(clk), .input_share0(d21_i21_s0), .input_share1(d21_i21_s1), .output_share0(d22_i21_s0), .output_share1(d22_i21_s1));
  reg_module u_reg_i22_d22 (.clk(clk), .input_share0(d21_i22_s0), .input_share1(d21_i22_s1), .output_share0(d22_i22_s0), .output_share1(d22_i22_s1));
  reg_module u_reg_i23_d22 (.clk(clk), .input_share0(d21_i23_s0), .input_share1(d21_i23_s1), .output_share0(d22_i23_s0), .output_share1(d22_i23_s1));
  reg_module u_reg_i24_d22 (.clk(clk), .input_share0(d21_i24_s0), .input_share1(d21_i24_s1), .output_share0(d22_i24_s0), .output_share1(d22_i24_s1));
  reg_module u_reg_i25_d22 (.clk(clk), .input_share0(d21_i25_s0), .input_share1(d21_i25_s1), .output_share0(d22_i25_s0), .output_share1(d22_i25_s1));
  reg_module u_reg_i26_d22 (.clk(clk), .input_share0(d21_i26_s0), .input_share1(d21_i26_s1), .output_share0(d22_i26_s0), .output_share1(d22_i26_s1));
  reg_module u_reg_i27_d22 (.clk(clk), .input_share0(d21_i27_s0), .input_share1(d21_i27_s1), .output_share0(d22_i27_s0), .output_share1(d22_i27_s1));
  reg_module u_reg_i28_d22 (.clk(clk), .input_share0(d21_i28_s0), .input_share1(d21_i28_s1), .output_share0(d22_i28_s0), .output_share1(d22_i28_s1));
  reg_module u_reg_i29_d22 (.clk(clk), .input_share0(d21_i29_s0), .input_share1(d21_i29_s1), .output_share0(d22_i29_s0), .output_share1(d22_i29_s1));
  reg_module u_reg_i30_d22 (.clk(clk), .input_share0(d21_i30_s0), .input_share1(d21_i30_s1), .output_share0(d22_i30_s0), .output_share1(d22_i30_s1));
  reg_module u_reg_t0_22_d22 (.clk(clk), .input_share0(d21_t0_22_s0), .input_share1(d21_t0_22_s1), .output_share0(d22_t0_22_s0), .output_share1(d22_t0_22_s1));
  reg_module u_reg_t0_23_d22 (.clk(clk), .input_share0(d21_t0_23_s0), .input_share1(d21_t0_23_s1), .output_share0(d22_t0_23_s0), .output_share1(d22_t0_23_s1));
  reg_module u_reg_t0_24_d22 (.clk(clk), .input_share0(d21_t0_24_s0), .input_share1(d21_t0_24_s1), .output_share0(d22_t0_24_s0), .output_share1(d22_t0_24_s1));
  reg_module u_reg_t0_25_d22 (.clk(clk), .input_share0(d21_t0_25_s0), .input_share1(d21_t0_25_s1), .output_share0(d22_t0_25_s0), .output_share1(d22_t0_25_s1));
  reg_module u_reg_t0_26_d22 (.clk(clk), .input_share0(d21_t0_26_s0), .input_share1(d21_t0_26_s1), .output_share0(d22_t0_26_s0), .output_share1(d22_t0_26_s1));
  reg_module u_reg_t0_27_d22 (.clk(clk), .input_share0(d21_t0_27_s0), .input_share1(d21_t0_27_s1), .output_share0(d22_t0_27_s0), .output_share1(d22_t0_27_s1));
  reg_module u_reg_t0_28_d22 (.clk(clk), .input_share0(d21_t0_28_s0), .input_share1(d21_t0_28_s1), .output_share0(d22_t0_28_s0), .output_share1(d22_t0_28_s1));
  reg_module u_reg_t0_29_d22 (.clk(clk), .input_share0(d21_t0_29_s0), .input_share1(d21_t0_29_s1), .output_share0(d22_t0_29_s0), .output_share1(d22_t0_29_s1));
  reg_module u_reg_t0_30_d22 (.clk(clk), .input_share0(d21_t0_30_s0), .input_share1(d21_t0_30_s1), .output_share0(d22_t0_30_s0), .output_share1(d22_t0_30_s1));
  reg_module u_reg_t0_31_d22 (.clk(clk), .input_share0(d21_t0_31_s0), .input_share1(d21_t0_31_s1), .output_share0(d22_t0_31_s0), .output_share1(d22_t0_31_s1));
  xor_module u_xor_c22_d22 (.x_share0(d22_i21_s0), .x_share1(d22_i21_s1), .y_share0(d22_t2_21_s0), .y_share1(d22_t2_21_s1), .z_share0(d22_c22_s0), .z_share1(d22_c22_s1));
  xor_module u_xor_o22_d22 (.x_share0(d22_t0_22_s0), .x_share1(d22_t0_22_s1), .y_share0(d22_c22_s0), .y_share1(d22_c22_s1), .z_share0(d22_o22_s0), .z_share1(d22_o22_s1));
  xor_module u_xor_t1_22_d22 (.x_share0(d22_i22_s0), .x_share1(d22_i22_s1), .y_share0(d22_c22_s0), .y_share1(d22_c22_s1), .z_share0(d22_t1_22_s0), .z_share1(d22_t1_22_s1));
  and_module u_and_t2_21_d22 (.clk(clk), .x_share0(d21_t0_21_s0), .x_share1(d21_t0_21_s1), .y_share0(d21_t1_21_s0), .y_share1(d21_t1_21_s1), .rand(r_t2_21), .z_share0(d22_t2_21_s0), .z_share1(d22_t2_21_s1));
  assign r_t2_21 = stage22_share0[1];
  reg_module u_reg_i22_d23 (.clk(clk), .input_share0(d22_i22_s0), .input_share1(d22_i22_s1), .output_share0(d23_i22_s0), .output_share1(d23_i22_s1));
  reg_module u_reg_i23_d23 (.clk(clk), .input_share0(d22_i23_s0), .input_share1(d22_i23_s1), .output_share0(d23_i23_s0), .output_share1(d23_i23_s1));
  reg_module u_reg_i24_d23 (.clk(clk), .input_share0(d22_i24_s0), .input_share1(d22_i24_s1), .output_share0(d23_i24_s0), .output_share1(d23_i24_s1));
  reg_module u_reg_i25_d23 (.clk(clk), .input_share0(d22_i25_s0), .input_share1(d22_i25_s1), .output_share0(d23_i25_s0), .output_share1(d23_i25_s1));
  reg_module u_reg_i26_d23 (.clk(clk), .input_share0(d22_i26_s0), .input_share1(d22_i26_s1), .output_share0(d23_i26_s0), .output_share1(d23_i26_s1));
  reg_module u_reg_i27_d23 (.clk(clk), .input_share0(d22_i27_s0), .input_share1(d22_i27_s1), .output_share0(d23_i27_s0), .output_share1(d23_i27_s1));
  reg_module u_reg_i28_d23 (.clk(clk), .input_share0(d22_i28_s0), .input_share1(d22_i28_s1), .output_share0(d23_i28_s0), .output_share1(d23_i28_s1));
  reg_module u_reg_i29_d23 (.clk(clk), .input_share0(d22_i29_s0), .input_share1(d22_i29_s1), .output_share0(d23_i29_s0), .output_share1(d23_i29_s1));
  reg_module u_reg_i30_d23 (.clk(clk), .input_share0(d22_i30_s0), .input_share1(d22_i30_s1), .output_share0(d23_i30_s0), .output_share1(d23_i30_s1));
  reg_module u_reg_t0_23_d23 (.clk(clk), .input_share0(d22_t0_23_s0), .input_share1(d22_t0_23_s1), .output_share0(d23_t0_23_s0), .output_share1(d23_t0_23_s1));
  reg_module u_reg_t0_24_d23 (.clk(clk), .input_share0(d22_t0_24_s0), .input_share1(d22_t0_24_s1), .output_share0(d23_t0_24_s0), .output_share1(d23_t0_24_s1));
  reg_module u_reg_t0_25_d23 (.clk(clk), .input_share0(d22_t0_25_s0), .input_share1(d22_t0_25_s1), .output_share0(d23_t0_25_s0), .output_share1(d23_t0_25_s1));
  reg_module u_reg_t0_26_d23 (.clk(clk), .input_share0(d22_t0_26_s0), .input_share1(d22_t0_26_s1), .output_share0(d23_t0_26_s0), .output_share1(d23_t0_26_s1));
  reg_module u_reg_t0_27_d23 (.clk(clk), .input_share0(d22_t0_27_s0), .input_share1(d22_t0_27_s1), .output_share0(d23_t0_27_s0), .output_share1(d23_t0_27_s1));
  reg_module u_reg_t0_28_d23 (.clk(clk), .input_share0(d22_t0_28_s0), .input_share1(d22_t0_28_s1), .output_share0(d23_t0_28_s0), .output_share1(d23_t0_28_s1));
  reg_module u_reg_t0_29_d23 (.clk(clk), .input_share0(d22_t0_29_s0), .input_share1(d22_t0_29_s1), .output_share0(d23_t0_29_s0), .output_share1(d23_t0_29_s1));
  reg_module u_reg_t0_30_d23 (.clk(clk), .input_share0(d22_t0_30_s0), .input_share1(d22_t0_30_s1), .output_share0(d23_t0_30_s0), .output_share1(d23_t0_30_s1));
  reg_module u_reg_t0_31_d23 (.clk(clk), .input_share0(d22_t0_31_s0), .input_share1(d22_t0_31_s1), .output_share0(d23_t0_31_s0), .output_share1(d23_t0_31_s1));
  xor_module u_xor_c23_d23 (.x_share0(d23_i22_s0), .x_share1(d23_i22_s1), .y_share0(d23_t2_22_s0), .y_share1(d23_t2_22_s1), .z_share0(d23_c23_s0), .z_share1(d23_c23_s1));
  xor_module u_xor_o23_d23 (.x_share0(d23_t0_23_s0), .x_share1(d23_t0_23_s1), .y_share0(d23_c23_s0), .y_share1(d23_c23_s1), .z_share0(d23_o23_s0), .z_share1(d23_o23_s1));
  xor_module u_xor_t1_23_d23 (.x_share0(d23_i23_s0), .x_share1(d23_i23_s1), .y_share0(d23_c23_s0), .y_share1(d23_c23_s1), .z_share0(d23_t1_23_s0), .z_share1(d23_t1_23_s1));
  and_module u_and_t2_22_d23 (.clk(clk), .x_share0(d22_t0_22_s0), .x_share1(d22_t0_22_s1), .y_share0(d22_t1_22_s0), .y_share1(d22_t1_22_s1), .rand(r_t2_22), .z_share0(d23_t2_22_s0), .z_share1(d23_t2_22_s1));
  assign r_t2_22 = stage23_share0[2];
  reg_module u_reg_i23_d24 (.clk(clk), .input_share0(d23_i23_s0), .input_share1(d23_i23_s1), .output_share0(d24_i23_s0), .output_share1(d24_i23_s1));
  reg_module u_reg_i24_d24 (.clk(clk), .input_share0(d23_i24_s0), .input_share1(d23_i24_s1), .output_share0(d24_i24_s0), .output_share1(d24_i24_s1));
  reg_module u_reg_i25_d24 (.clk(clk), .input_share0(d23_i25_s0), .input_share1(d23_i25_s1), .output_share0(d24_i25_s0), .output_share1(d24_i25_s1));
  reg_module u_reg_i26_d24 (.clk(clk), .input_share0(d23_i26_s0), .input_share1(d23_i26_s1), .output_share0(d24_i26_s0), .output_share1(d24_i26_s1));
  reg_module u_reg_i27_d24 (.clk(clk), .input_share0(d23_i27_s0), .input_share1(d23_i27_s1), .output_share0(d24_i27_s0), .output_share1(d24_i27_s1));
  reg_module u_reg_i28_d24 (.clk(clk), .input_share0(d23_i28_s0), .input_share1(d23_i28_s1), .output_share0(d24_i28_s0), .output_share1(d24_i28_s1));
  reg_module u_reg_i29_d24 (.clk(clk), .input_share0(d23_i29_s0), .input_share1(d23_i29_s1), .output_share0(d24_i29_s0), .output_share1(d24_i29_s1));
  reg_module u_reg_i30_d24 (.clk(clk), .input_share0(d23_i30_s0), .input_share1(d23_i30_s1), .output_share0(d24_i30_s0), .output_share1(d24_i30_s1));
  reg_module u_reg_t0_24_d24 (.clk(clk), .input_share0(d23_t0_24_s0), .input_share1(d23_t0_24_s1), .output_share0(d24_t0_24_s0), .output_share1(d24_t0_24_s1));
  reg_module u_reg_t0_25_d24 (.clk(clk), .input_share0(d23_t0_25_s0), .input_share1(d23_t0_25_s1), .output_share0(d24_t0_25_s0), .output_share1(d24_t0_25_s1));
  reg_module u_reg_t0_26_d24 (.clk(clk), .input_share0(d23_t0_26_s0), .input_share1(d23_t0_26_s1), .output_share0(d24_t0_26_s0), .output_share1(d24_t0_26_s1));
  reg_module u_reg_t0_27_d24 (.clk(clk), .input_share0(d23_t0_27_s0), .input_share1(d23_t0_27_s1), .output_share0(d24_t0_27_s0), .output_share1(d24_t0_27_s1));
  reg_module u_reg_t0_28_d24 (.clk(clk), .input_share0(d23_t0_28_s0), .input_share1(d23_t0_28_s1), .output_share0(d24_t0_28_s0), .output_share1(d24_t0_28_s1));
  reg_module u_reg_t0_29_d24 (.clk(clk), .input_share0(d23_t0_29_s0), .input_share1(d23_t0_29_s1), .output_share0(d24_t0_29_s0), .output_share1(d24_t0_29_s1));
  reg_module u_reg_t0_30_d24 (.clk(clk), .input_share0(d23_t0_30_s0), .input_share1(d23_t0_30_s1), .output_share0(d24_t0_30_s0), .output_share1(d24_t0_30_s1));
  reg_module u_reg_t0_31_d24 (.clk(clk), .input_share0(d23_t0_31_s0), .input_share1(d23_t0_31_s1), .output_share0(d24_t0_31_s0), .output_share1(d24_t0_31_s1));
  xor_module u_xor_c24_d24 (.x_share0(d24_i23_s0), .x_share1(d24_i23_s1), .y_share0(d24_t2_23_s0), .y_share1(d24_t2_23_s1), .z_share0(d24_c24_s0), .z_share1(d24_c24_s1));
  xor_module u_xor_o24_d24 (.x_share0(d24_t0_24_s0), .x_share1(d24_t0_24_s1), .y_share0(d24_c24_s0), .y_share1(d24_c24_s1), .z_share0(d24_o24_s0), .z_share1(d24_o24_s1));
  xor_module u_xor_t1_24_d24 (.x_share0(d24_i24_s0), .x_share1(d24_i24_s1), .y_share0(d24_c24_s0), .y_share1(d24_c24_s1), .z_share0(d24_t1_24_s0), .z_share1(d24_t1_24_s1));
  and_module u_and_t2_23_d24 (.clk(clk), .x_share0(d23_t0_23_s0), .x_share1(d23_t0_23_s1), .y_share0(d23_t1_23_s0), .y_share1(d23_t1_23_s1), .rand(r_t2_23), .z_share0(d24_t2_23_s0), .z_share1(d24_t2_23_s1));
  assign r_t2_23 = stage24_share0[0];
  reg_module u_reg_i24_d25 (.clk(clk), .input_share0(d24_i24_s0), .input_share1(d24_i24_s1), .output_share0(d25_i24_s0), .output_share1(d25_i24_s1));
  reg_module u_reg_i25_d25 (.clk(clk), .input_share0(d24_i25_s0), .input_share1(d24_i25_s1), .output_share0(d25_i25_s0), .output_share1(d25_i25_s1));
  reg_module u_reg_i26_d25 (.clk(clk), .input_share0(d24_i26_s0), .input_share1(d24_i26_s1), .output_share0(d25_i26_s0), .output_share1(d25_i26_s1));
  reg_module u_reg_i27_d25 (.clk(clk), .input_share0(d24_i27_s0), .input_share1(d24_i27_s1), .output_share0(d25_i27_s0), .output_share1(d25_i27_s1));
  reg_module u_reg_i28_d25 (.clk(clk), .input_share0(d24_i28_s0), .input_share1(d24_i28_s1), .output_share0(d25_i28_s0), .output_share1(d25_i28_s1));
  reg_module u_reg_i29_d25 (.clk(clk), .input_share0(d24_i29_s0), .input_share1(d24_i29_s1), .output_share0(d25_i29_s0), .output_share1(d25_i29_s1));
  reg_module u_reg_i30_d25 (.clk(clk), .input_share0(d24_i30_s0), .input_share1(d24_i30_s1), .output_share0(d25_i30_s0), .output_share1(d25_i30_s1));
  reg_module u_reg_t0_25_d25 (.clk(clk), .input_share0(d24_t0_25_s0), .input_share1(d24_t0_25_s1), .output_share0(d25_t0_25_s0), .output_share1(d25_t0_25_s1));
  reg_module u_reg_t0_26_d25 (.clk(clk), .input_share0(d24_t0_26_s0), .input_share1(d24_t0_26_s1), .output_share0(d25_t0_26_s0), .output_share1(d25_t0_26_s1));
  reg_module u_reg_t0_27_d25 (.clk(clk), .input_share0(d24_t0_27_s0), .input_share1(d24_t0_27_s1), .output_share0(d25_t0_27_s0), .output_share1(d25_t0_27_s1));
  reg_module u_reg_t0_28_d25 (.clk(clk), .input_share0(d24_t0_28_s0), .input_share1(d24_t0_28_s1), .output_share0(d25_t0_28_s0), .output_share1(d25_t0_28_s1));
  reg_module u_reg_t0_29_d25 (.clk(clk), .input_share0(d24_t0_29_s0), .input_share1(d24_t0_29_s1), .output_share0(d25_t0_29_s0), .output_share1(d25_t0_29_s1));
  reg_module u_reg_t0_30_d25 (.clk(clk), .input_share0(d24_t0_30_s0), .input_share1(d24_t0_30_s1), .output_share0(d25_t0_30_s0), .output_share1(d25_t0_30_s1));
  reg_module u_reg_t0_31_d25 (.clk(clk), .input_share0(d24_t0_31_s0), .input_share1(d24_t0_31_s1), .output_share0(d25_t0_31_s0), .output_share1(d25_t0_31_s1));
  xor_module u_xor_c25_d25 (.x_share0(d25_i24_s0), .x_share1(d25_i24_s1), .y_share0(d25_t2_24_s0), .y_share1(d25_t2_24_s1), .z_share0(d25_c25_s0), .z_share1(d25_c25_s1));
  xor_module u_xor_o25_d25 (.x_share0(d25_t0_25_s0), .x_share1(d25_t0_25_s1), .y_share0(d25_c25_s0), .y_share1(d25_c25_s1), .z_share0(d25_o25_s0), .z_share1(d25_o25_s1));
  xor_module u_xor_t1_25_d25 (.x_share0(d25_i25_s0), .x_share1(d25_i25_s1), .y_share0(d25_c25_s0), .y_share1(d25_c25_s1), .z_share0(d25_t1_25_s0), .z_share1(d25_t1_25_s1));
  and_module u_and_t2_24_d25 (.clk(clk), .x_share0(d24_t0_24_s0), .x_share1(d24_t0_24_s1), .y_share0(d24_t1_24_s0), .y_share1(d24_t1_24_s1), .rand(r_t2_24), .z_share0(d25_t2_24_s0), .z_share1(d25_t2_24_s1));
  assign r_t2_24 = stage25_share0[1];
  reg_module u_reg_i25_d26 (.clk(clk), .input_share0(d25_i25_s0), .input_share1(d25_i25_s1), .output_share0(d26_i25_s0), .output_share1(d26_i25_s1));
  reg_module u_reg_i26_d26 (.clk(clk), .input_share0(d25_i26_s0), .input_share1(d25_i26_s1), .output_share0(d26_i26_s0), .output_share1(d26_i26_s1));
  reg_module u_reg_i27_d26 (.clk(clk), .input_share0(d25_i27_s0), .input_share1(d25_i27_s1), .output_share0(d26_i27_s0), .output_share1(d26_i27_s1));
  reg_module u_reg_i28_d26 (.clk(clk), .input_share0(d25_i28_s0), .input_share1(d25_i28_s1), .output_share0(d26_i28_s0), .output_share1(d26_i28_s1));
  reg_module u_reg_i29_d26 (.clk(clk), .input_share0(d25_i29_s0), .input_share1(d25_i29_s1), .output_share0(d26_i29_s0), .output_share1(d26_i29_s1));
  reg_module u_reg_i30_d26 (.clk(clk), .input_share0(d25_i30_s0), .input_share1(d25_i30_s1), .output_share0(d26_i30_s0), .output_share1(d26_i30_s1));
  reg_module u_reg_t0_26_d26 (.clk(clk), .input_share0(d25_t0_26_s0), .input_share1(d25_t0_26_s1), .output_share0(d26_t0_26_s0), .output_share1(d26_t0_26_s1));
  reg_module u_reg_t0_27_d26 (.clk(clk), .input_share0(d25_t0_27_s0), .input_share1(d25_t0_27_s1), .output_share0(d26_t0_27_s0), .output_share1(d26_t0_27_s1));
  reg_module u_reg_t0_28_d26 (.clk(clk), .input_share0(d25_t0_28_s0), .input_share1(d25_t0_28_s1), .output_share0(d26_t0_28_s0), .output_share1(d26_t0_28_s1));
  reg_module u_reg_t0_29_d26 (.clk(clk), .input_share0(d25_t0_29_s0), .input_share1(d25_t0_29_s1), .output_share0(d26_t0_29_s0), .output_share1(d26_t0_29_s1));
  reg_module u_reg_t0_30_d26 (.clk(clk), .input_share0(d25_t0_30_s0), .input_share1(d25_t0_30_s1), .output_share0(d26_t0_30_s0), .output_share1(d26_t0_30_s1));
  reg_module u_reg_t0_31_d26 (.clk(clk), .input_share0(d25_t0_31_s0), .input_share1(d25_t0_31_s1), .output_share0(d26_t0_31_s0), .output_share1(d26_t0_31_s1));
  xor_module u_xor_c26_d26 (.x_share0(d26_i25_s0), .x_share1(d26_i25_s1), .y_share0(d26_t2_25_s0), .y_share1(d26_t2_25_s1), .z_share0(d26_c26_s0), .z_share1(d26_c26_s1));
  xor_module u_xor_o26_d26 (.x_share0(d26_t0_26_s0), .x_share1(d26_t0_26_s1), .y_share0(d26_c26_s0), .y_share1(d26_c26_s1), .z_share0(d26_o26_s0), .z_share1(d26_o26_s1));
  xor_module u_xor_t1_26_d26 (.x_share0(d26_i26_s0), .x_share1(d26_i26_s1), .y_share0(d26_c26_s0), .y_share1(d26_c26_s1), .z_share0(d26_t1_26_s0), .z_share1(d26_t1_26_s1));
  and_module u_and_t2_25_d26 (.clk(clk), .x_share0(d25_t0_25_s0), .x_share1(d25_t0_25_s1), .y_share0(d25_t1_25_s0), .y_share1(d25_t1_25_s1), .rand(r_t2_25), .z_share0(d26_t2_25_s0), .z_share1(d26_t2_25_s1));
  assign r_t2_25 = stage26_share0[2];
  reg_module u_reg_i26_d27 (.clk(clk), .input_share0(d26_i26_s0), .input_share1(d26_i26_s1), .output_share0(d27_i26_s0), .output_share1(d27_i26_s1));
  reg_module u_reg_i27_d27 (.clk(clk), .input_share0(d26_i27_s0), .input_share1(d26_i27_s1), .output_share0(d27_i27_s0), .output_share1(d27_i27_s1));
  reg_module u_reg_i28_d27 (.clk(clk), .input_share0(d26_i28_s0), .input_share1(d26_i28_s1), .output_share0(d27_i28_s0), .output_share1(d27_i28_s1));
  reg_module u_reg_i29_d27 (.clk(clk), .input_share0(d26_i29_s0), .input_share1(d26_i29_s1), .output_share0(d27_i29_s0), .output_share1(d27_i29_s1));
  reg_module u_reg_i30_d27 (.clk(clk), .input_share0(d26_i30_s0), .input_share1(d26_i30_s1), .output_share0(d27_i30_s0), .output_share1(d27_i30_s1));
  reg_module u_reg_t0_27_d27 (.clk(clk), .input_share0(d26_t0_27_s0), .input_share1(d26_t0_27_s1), .output_share0(d27_t0_27_s0), .output_share1(d27_t0_27_s1));
  reg_module u_reg_t0_28_d27 (.clk(clk), .input_share0(d26_t0_28_s0), .input_share1(d26_t0_28_s1), .output_share0(d27_t0_28_s0), .output_share1(d27_t0_28_s1));
  reg_module u_reg_t0_29_d27 (.clk(clk), .input_share0(d26_t0_29_s0), .input_share1(d26_t0_29_s1), .output_share0(d27_t0_29_s0), .output_share1(d27_t0_29_s1));
  reg_module u_reg_t0_30_d27 (.clk(clk), .input_share0(d26_t0_30_s0), .input_share1(d26_t0_30_s1), .output_share0(d27_t0_30_s0), .output_share1(d27_t0_30_s1));
  reg_module u_reg_t0_31_d27 (.clk(clk), .input_share0(d26_t0_31_s0), .input_share1(d26_t0_31_s1), .output_share0(d27_t0_31_s0), .output_share1(d27_t0_31_s1));
  xor_module u_xor_c27_d27 (.x_share0(d27_i26_s0), .x_share1(d27_i26_s1), .y_share0(d27_t2_26_s0), .y_share1(d27_t2_26_s1), .z_share0(d27_c27_s0), .z_share1(d27_c27_s1));
  xor_module u_xor_o27_d27 (.x_share0(d27_t0_27_s0), .x_share1(d27_t0_27_s1), .y_share0(d27_c27_s0), .y_share1(d27_c27_s1), .z_share0(d27_o27_s0), .z_share1(d27_o27_s1));
  xor_module u_xor_t1_27_d27 (.x_share0(d27_i27_s0), .x_share1(d27_i27_s1), .y_share0(d27_c27_s0), .y_share1(d27_c27_s1), .z_share0(d27_t1_27_s0), .z_share1(d27_t1_27_s1));
  and_module u_and_t2_26_d27 (.clk(clk), .x_share0(d26_t0_26_s0), .x_share1(d26_t0_26_s1), .y_share0(d26_t1_26_s0), .y_share1(d26_t1_26_s1), .rand(r_t2_26), .z_share0(d27_t2_26_s0), .z_share1(d27_t2_26_s1));
  assign r_t2_26 = stage27_share0[0];
  reg_module u_reg_i27_d28 (.clk(clk), .input_share0(d27_i27_s0), .input_share1(d27_i27_s1), .output_share0(d28_i27_s0), .output_share1(d28_i27_s1));
  reg_module u_reg_i28_d28 (.clk(clk), .input_share0(d27_i28_s0), .input_share1(d27_i28_s1), .output_share0(d28_i28_s0), .output_share1(d28_i28_s1));
  reg_module u_reg_i29_d28 (.clk(clk), .input_share0(d27_i29_s0), .input_share1(d27_i29_s1), .output_share0(d28_i29_s0), .output_share1(d28_i29_s1));
  reg_module u_reg_i30_d28 (.clk(clk), .input_share0(d27_i30_s0), .input_share1(d27_i30_s1), .output_share0(d28_i30_s0), .output_share1(d28_i30_s1));
  reg_module u_reg_t0_28_d28 (.clk(clk), .input_share0(d27_t0_28_s0), .input_share1(d27_t0_28_s1), .output_share0(d28_t0_28_s0), .output_share1(d28_t0_28_s1));
  reg_module u_reg_t0_29_d28 (.clk(clk), .input_share0(d27_t0_29_s0), .input_share1(d27_t0_29_s1), .output_share0(d28_t0_29_s0), .output_share1(d28_t0_29_s1));
  reg_module u_reg_t0_30_d28 (.clk(clk), .input_share0(d27_t0_30_s0), .input_share1(d27_t0_30_s1), .output_share0(d28_t0_30_s0), .output_share1(d28_t0_30_s1));
  reg_module u_reg_t0_31_d28 (.clk(clk), .input_share0(d27_t0_31_s0), .input_share1(d27_t0_31_s1), .output_share0(d28_t0_31_s0), .output_share1(d28_t0_31_s1));
  xor_module u_xor_c28_d28 (.x_share0(d28_i27_s0), .x_share1(d28_i27_s1), .y_share0(d28_t2_27_s0), .y_share1(d28_t2_27_s1), .z_share0(d28_c28_s0), .z_share1(d28_c28_s1));
  xor_module u_xor_o28_d28 (.x_share0(d28_t0_28_s0), .x_share1(d28_t0_28_s1), .y_share0(d28_c28_s0), .y_share1(d28_c28_s1), .z_share0(d28_o28_s0), .z_share1(d28_o28_s1));
  xor_module u_xor_t1_28_d28 (.x_share0(d28_i28_s0), .x_share1(d28_i28_s1), .y_share0(d28_c28_s0), .y_share1(d28_c28_s1), .z_share0(d28_t1_28_s0), .z_share1(d28_t1_28_s1));
  and_module u_and_t2_27_d28 (.clk(clk), .x_share0(d27_t0_27_s0), .x_share1(d27_t0_27_s1), .y_share0(d27_t1_27_s0), .y_share1(d27_t1_27_s1), .rand(r_t2_27), .z_share0(d28_t2_27_s0), .z_share1(d28_t2_27_s1));
  assign r_t2_27 = stage28_share0[1];
  reg_module u_reg_i28_d29 (.clk(clk), .input_share0(d28_i28_s0), .input_share1(d28_i28_s1), .output_share0(d29_i28_s0), .output_share1(d29_i28_s1));
  reg_module u_reg_i29_d29 (.clk(clk), .input_share0(d28_i29_s0), .input_share1(d28_i29_s1), .output_share0(d29_i29_s0), .output_share1(d29_i29_s1));
  reg_module u_reg_i30_d29 (.clk(clk), .input_share0(d28_i30_s0), .input_share1(d28_i30_s1), .output_share0(d29_i30_s0), .output_share1(d29_i30_s1));
  reg_module u_reg_t0_29_d29 (.clk(clk), .input_share0(d28_t0_29_s0), .input_share1(d28_t0_29_s1), .output_share0(d29_t0_29_s0), .output_share1(d29_t0_29_s1));
  reg_module u_reg_t0_30_d29 (.clk(clk), .input_share0(d28_t0_30_s0), .input_share1(d28_t0_30_s1), .output_share0(d29_t0_30_s0), .output_share1(d29_t0_30_s1));
  reg_module u_reg_t0_31_d29 (.clk(clk), .input_share0(d28_t0_31_s0), .input_share1(d28_t0_31_s1), .output_share0(d29_t0_31_s0), .output_share1(d29_t0_31_s1));
  xor_module u_xor_c29_d29 (.x_share0(d29_i28_s0), .x_share1(d29_i28_s1), .y_share0(d29_t2_28_s0), .y_share1(d29_t2_28_s1), .z_share0(d29_c29_s0), .z_share1(d29_c29_s1));
  xor_module u_xor_o29_d29 (.x_share0(d29_t0_29_s0), .x_share1(d29_t0_29_s1), .y_share0(d29_c29_s0), .y_share1(d29_c29_s1), .z_share0(d29_o29_s0), .z_share1(d29_o29_s1));
  xor_module u_xor_t1_29_d29 (.x_share0(d29_i29_s0), .x_share1(d29_i29_s1), .y_share0(d29_c29_s0), .y_share1(d29_c29_s1), .z_share0(d29_t1_29_s0), .z_share1(d29_t1_29_s1));
  and_module u_and_t2_28_d29 (.clk(clk), .x_share0(d28_t0_28_s0), .x_share1(d28_t0_28_s1), .y_share0(d28_t1_28_s0), .y_share1(d28_t1_28_s1), .rand(r_t2_28), .z_share0(d29_t2_28_s0), .z_share1(d29_t2_28_s1));
  assign r_t2_28 = stage29_share0[2];
  reg_module u_reg_i29_d30 (.clk(clk), .input_share0(d29_i29_s0), .input_share1(d29_i29_s1), .output_share0(d30_i29_s0), .output_share1(d30_i29_s1));
  reg_module u_reg_i30_d30 (.clk(clk), .input_share0(d29_i30_s0), .input_share1(d29_i30_s1), .output_share0(d30_i30_s0), .output_share1(d30_i30_s1));
  reg_module u_reg_t0_30_d30 (.clk(clk), .input_share0(d29_t0_30_s0), .input_share1(d29_t0_30_s1), .output_share0(d30_t0_30_s0), .output_share1(d30_t0_30_s1));
  reg_module u_reg_t0_31_d30 (.clk(clk), .input_share0(d29_t0_31_s0), .input_share1(d29_t0_31_s1), .output_share0(d30_t0_31_s0), .output_share1(d30_t0_31_s1));
  xor_module u_xor_c30_d30 (.x_share0(d30_i29_s0), .x_share1(d30_i29_s1), .y_share0(d30_t2_29_s0), .y_share1(d30_t2_29_s1), .z_share0(d30_c30_s0), .z_share1(d30_c30_s1));
  xor_module u_xor_o30_d30 (.x_share0(d30_t0_30_s0), .x_share1(d30_t0_30_s1), .y_share0(d30_c30_s0), .y_share1(d30_c30_s1), .z_share0(d30_o30_s0), .z_share1(d30_o30_s1));
  xor_module u_xor_t1_30_d30 (.x_share0(d30_i30_s0), .x_share1(d30_i30_s1), .y_share0(d30_c30_s0), .y_share1(d30_c30_s1), .z_share0(d30_t1_30_s0), .z_share1(d30_t1_30_s1));
  and_module u_and_t2_29_d30 (.clk(clk), .x_share0(d29_t0_29_s0), .x_share1(d29_t0_29_s1), .y_share0(d29_t1_29_s0), .y_share1(d29_t1_29_s1), .rand(r_t2_29), .z_share0(d30_t2_29_s0), .z_share1(d30_t2_29_s1));
  assign r_t2_29 = stage30_share0[0];
  reg_module u_reg_i30_d31 (.clk(clk), .input_share0(d30_i30_s0), .input_share1(d30_i30_s1), .output_share0(d31_i30_s0), .output_share1(d31_i30_s1));
  reg_module u_reg_t0_31_d31 (.clk(clk), .input_share0(d30_t0_31_s0), .input_share1(d30_t0_31_s1), .output_share0(d31_t0_31_s0), .output_share1(d31_t0_31_s1));
  xor_module u_xor_c31_d31 (.x_share0(d31_i30_s0), .x_share1(d31_i30_s1), .y_share0(d31_t2_30_s0), .y_share1(d31_t2_30_s1), .z_share0(d31_c31_s0), .z_share1(d31_c31_s1));
  xor_module u_xor_o31_d31 (.x_share0(d31_t0_31_s0), .x_share1(d31_t0_31_s1), .y_share0(d31_c31_s0), .y_share1(d31_c31_s1), .z_share0(d31_o31_s0), .z_share1(d31_o31_s1));
  and_module u_and_t2_30_d31 (.clk(clk), .x_share0(d30_t0_30_s0), .x_share1(d30_t0_30_s1), .y_share0(d30_t1_30_s0), .y_share1(d30_t1_30_s1), .rand(r_t2_30), .z_share0(d31_t2_30_s0), .z_share1(d31_t2_30_s1));
  assign r_t2_30 = stage31_share0[1];

  // Output assignments
  assign o_share0[0] = d0_o0_s0;
  assign o_share1[0] = d0_o0_s1;
  assign o_share0[1] = d1_o1_s0;
  assign o_share1[1] = d1_o1_s1;
  assign o_share0[2] = d2_o2_s0;
  assign o_share1[2] = d2_o2_s1;
  assign o_share0[3] = d3_o3_s0;
  assign o_share1[3] = d3_o3_s1;
  assign o_share0[4] = d4_o4_s0;
  assign o_share1[4] = d4_o4_s1;
  assign o_share0[5] = d5_o5_s0;
  assign o_share1[5] = d5_o5_s1;
  assign o_share0[6] = d6_o6_s0;
  assign o_share1[6] = d6_o6_s1;
  assign o_share0[7] = d7_o7_s0;
  assign o_share1[7] = d7_o7_s1;
  assign o_share0[8] = d8_o8_s0;
  assign o_share1[8] = d8_o8_s1;
  assign o_share0[9] = d9_o9_s0;
  assign o_share1[9] = d9_o9_s1;
  assign o_share0[10] = d10_o10_s0;
  assign o_share1[10] = d10_o10_s1;
  assign o_share0[11] = d11_o11_s0;
  assign o_share1[11] = d11_o11_s1;
  assign o_share0[12] = d12_o12_s0;
  assign o_share1[12] = d12_o12_s1;
  assign o_share0[13] = d13_o13_s0;
  assign o_share1[13] = d13_o13_s1;
  assign o_share0[14] = d14_o14_s0;
  assign o_share1[14] = d14_o14_s1;
  assign o_share0[15] = d15_o15_s0;
  assign o_share1[15] = d15_o15_s1;
  assign o_share0[16] = d16_o16_s0;
  assign o_share1[16] = d16_o16_s1;
  assign o_share0[17] = d17_o17_s0;
  assign o_share1[17] = d17_o17_s1;
  assign o_share0[18] = d18_o18_s0;
  assign o_share1[18] = d18_o18_s1;
  assign o_share0[19] = d19_o19_s0;
  assign o_share1[19] = d19_o19_s1;
  assign o_share0[20] = d20_o20_s0;
  assign o_share1[20] = d20_o20_s1;
  assign o_share0[21] = d21_o21_s0;
  assign o_share1[21] = d21_o21_s1;
  assign o_share0[22] = d22_o22_s0;
  assign o_share1[22] = d22_o22_s1;
  assign o_share0[23] = d23_o23_s0;
  assign o_share1[23] = d23_o23_s1;
  assign o_share0[24] = d24_o24_s0;
  assign o_share1[24] = d24_o24_s1;
  assign o_share0[25] = d25_o25_s0;
  assign o_share1[25] = d25_o25_s1;
  assign o_share0[26] = d26_o26_s0;
  assign o_share1[26] = d26_o26_s1;
  assign o_share0[27] = d27_o27_s0;
  assign o_share1[27] = d27_o27_s1;
  assign o_share0[28] = d28_o28_s0;
  assign o_share1[28] = d28_o28_s1;
  assign o_share0[29] = d29_o29_s0;
  assign o_share1[29] = d29_o29_s1;
  assign o_share0[30] = d30_o30_s0;
  assign o_share1[30] = d30_o30_s1;
  assign o_share0[31] = d31_o31_s0;
  assign o_share1[31] = d31_o31_s1;

endmodule
