`timescale 1ns / 1ps


module KSmod_32_latency_5 (
  input           clk,
  input  [63:0] share0_in,
  input  [63:0] share1_in,
  input  [26:0] rand_bit_share0,
  input  [26:0] rand_bit_share1,
  output [31:0] o_share0,
  output [31:0] o_share1
);

  // Randomness pipeline
  // depth-1 ANDs use rand_bit_share0 directly; deeper ones use these
  wire   [26:0] stage2_share0, stage3_share0, stage4_share0, stage5_share0, stage6_share0;

  reg_27bits rand_stage1 (.clk(clk), .input_share0(rand_bit_share0), .output_share0(stage2_share0));
  reg_27bits rand_stage2 (.clk(clk), .input_share0(stage2_share0), .output_share0(stage3_share0));
  reg_27bits rand_stage3 (.clk(clk), .input_share0(stage3_share0), .output_share0(stage4_share0));
  reg_27bits rand_stage4 (.clk(clk), .input_share0(stage4_share0), .output_share0(stage5_share0));
  reg_27bits rand_stage5 (.clk(clk), .input_share0(stage5_share0), .output_share0(stage6_share0));

  xor_module u_xor_P0_1_d0 (.x_share0(share0_in[1]), .x_share1(share1_in[1]), .y_share0(share0_in[33]), .y_share1(share1_in[33]), .z_share0(d0_P0_1_s0), .z_share1(d0_P0_1_s1));
  xor_module u_xor_P0_10_d0 (.x_share0(share0_in[10]), .x_share1(share1_in[10]), .y_share0(share0_in[42]), .y_share1(share1_in[42]), .z_share0(d0_P0_10_s0), .z_share1(d0_P0_10_s1));
  xor_module u_xor_P0_11_d0 (.x_share0(share0_in[11]), .x_share1(share1_in[11]), .y_share0(share0_in[43]), .y_share1(share1_in[43]), .z_share0(d0_P0_11_s0), .z_share1(d0_P0_11_s1));
  xor_module u_xor_P0_12_d0 (.x_share0(share0_in[12]), .x_share1(share1_in[12]), .y_share0(share0_in[44]), .y_share1(share1_in[44]), .z_share0(d0_P0_12_s0), .z_share1(d0_P0_12_s1));
  xor_module u_xor_P0_13_d0 (.x_share0(share0_in[13]), .x_share1(share1_in[13]), .y_share0(share0_in[45]), .y_share1(share1_in[45]), .z_share0(d0_P0_13_s0), .z_share1(d0_P0_13_s1));
  xor_module u_xor_P0_14_d0 (.x_share0(share0_in[14]), .x_share1(share1_in[14]), .y_share0(share0_in[46]), .y_share1(share1_in[46]), .z_share0(d0_P0_14_s0), .z_share1(d0_P0_14_s1));
  xor_module u_xor_P0_15_d0 (.x_share0(share0_in[15]), .x_share1(share1_in[15]), .y_share0(share0_in[47]), .y_share1(share1_in[47]), .z_share0(d0_P0_15_s0), .z_share1(d0_P0_15_s1));
  xor_module u_xor_P0_16_d0 (.x_share0(share0_in[16]), .x_share1(share1_in[16]), .y_share0(share0_in[48]), .y_share1(share1_in[48]), .z_share0(d0_P0_16_s0), .z_share1(d0_P0_16_s1));
  xor_module u_xor_P0_17_d0 (.x_share0(share0_in[17]), .x_share1(share1_in[17]), .y_share0(share0_in[49]), .y_share1(share1_in[49]), .z_share0(d0_P0_17_s0), .z_share1(d0_P0_17_s1));
  xor_module u_xor_P0_18_d0 (.x_share0(share0_in[18]), .x_share1(share1_in[18]), .y_share0(share0_in[50]), .y_share1(share1_in[50]), .z_share0(d0_P0_18_s0), .z_share1(d0_P0_18_s1));
  xor_module u_xor_P0_19_d0 (.x_share0(share0_in[19]), .x_share1(share1_in[19]), .y_share0(share0_in[51]), .y_share1(share1_in[51]), .z_share0(d0_P0_19_s0), .z_share1(d0_P0_19_s1));
  xor_module u_xor_P0_2_d0 (.x_share0(share0_in[2]), .x_share1(share1_in[2]), .y_share0(share0_in[34]), .y_share1(share1_in[34]), .z_share0(d0_P0_2_s0), .z_share1(d0_P0_2_s1));
  xor_module u_xor_P0_20_d0 (.x_share0(share0_in[20]), .x_share1(share1_in[20]), .y_share0(share0_in[52]), .y_share1(share1_in[52]), .z_share0(d0_P0_20_s0), .z_share1(d0_P0_20_s1));
  xor_module u_xor_P0_21_d0 (.x_share0(share0_in[21]), .x_share1(share1_in[21]), .y_share0(share0_in[53]), .y_share1(share1_in[53]), .z_share0(d0_P0_21_s0), .z_share1(d0_P0_21_s1));
  xor_module u_xor_P0_22_d0 (.x_share0(share0_in[22]), .x_share1(share1_in[22]), .y_share0(share0_in[54]), .y_share1(share1_in[54]), .z_share0(d0_P0_22_s0), .z_share1(d0_P0_22_s1));
  xor_module u_xor_P0_23_d0 (.x_share0(share0_in[23]), .x_share1(share1_in[23]), .y_share0(share0_in[55]), .y_share1(share1_in[55]), .z_share0(d0_P0_23_s0), .z_share1(d0_P0_23_s1));
  xor_module u_xor_P0_24_d0 (.x_share0(share0_in[24]), .x_share1(share1_in[24]), .y_share0(share0_in[56]), .y_share1(share1_in[56]), .z_share0(d0_P0_24_s0), .z_share1(d0_P0_24_s1));
  xor_module u_xor_P0_25_d0 (.x_share0(share0_in[25]), .x_share1(share1_in[25]), .y_share0(share0_in[57]), .y_share1(share1_in[57]), .z_share0(d0_P0_25_s0), .z_share1(d0_P0_25_s1));
  xor_module u_xor_P0_26_d0 (.x_share0(share0_in[26]), .x_share1(share1_in[26]), .y_share0(share0_in[58]), .y_share1(share1_in[58]), .z_share0(d0_P0_26_s0), .z_share1(d0_P0_26_s1));
  xor_module u_xor_P0_27_d0 (.x_share0(share0_in[27]), .x_share1(share1_in[27]), .y_share0(share0_in[59]), .y_share1(share1_in[59]), .z_share0(d0_P0_27_s0), .z_share1(d0_P0_27_s1));
  xor_module u_xor_P0_28_d0 (.x_share0(share0_in[28]), .x_share1(share1_in[28]), .y_share0(share0_in[60]), .y_share1(share1_in[60]), .z_share0(d0_P0_28_s0), .z_share1(d0_P0_28_s1));
  xor_module u_xor_P0_29_d0 (.x_share0(share0_in[29]), .x_share1(share1_in[29]), .y_share0(share0_in[61]), .y_share1(share1_in[61]), .z_share0(d0_P0_29_s0), .z_share1(d0_P0_29_s1));
  xor_module u_xor_P0_3_d0 (.x_share0(share0_in[3]), .x_share1(share1_in[3]), .y_share0(share0_in[35]), .y_share1(share1_in[35]), .z_share0(d0_P0_3_s0), .z_share1(d0_P0_3_s1));
  xor_module u_xor_P0_30_d0 (.x_share0(share0_in[30]), .x_share1(share1_in[30]), .y_share0(share0_in[62]), .y_share1(share1_in[62]), .z_share0(d0_P0_30_s0), .z_share1(d0_P0_30_s1));
  xor_module u_xor_P0_31_d0 (.x_share0(share0_in[31]), .x_share1(share1_in[31]), .y_share0(share0_in[63]), .y_share1(share1_in[63]), .z_share0(d0_P0_31_s0), .z_share1(d0_P0_31_s1));
  xor_module u_xor_P0_4_d0 (.x_share0(share0_in[4]), .x_share1(share1_in[4]), .y_share0(share0_in[36]), .y_share1(share1_in[36]), .z_share0(d0_P0_4_s0), .z_share1(d0_P0_4_s1));
  xor_module u_xor_P0_5_d0 (.x_share0(share0_in[5]), .x_share1(share1_in[5]), .y_share0(share0_in[37]), .y_share1(share1_in[37]), .z_share0(d0_P0_5_s0), .z_share1(d0_P0_5_s1));
  xor_module u_xor_P0_6_d0 (.x_share0(share0_in[6]), .x_share1(share1_in[6]), .y_share0(share0_in[38]), .y_share1(share1_in[38]), .z_share0(d0_P0_6_s0), .z_share1(d0_P0_6_s1));
  xor_module u_xor_P0_7_d0 (.x_share0(share0_in[7]), .x_share1(share1_in[7]), .y_share0(share0_in[39]), .y_share1(share1_in[39]), .z_share0(d0_P0_7_s0), .z_share1(d0_P0_7_s1));
  xor_module u_xor_P0_8_d0 (.x_share0(share0_in[8]), .x_share1(share1_in[8]), .y_share0(share0_in[40]), .y_share1(share1_in[40]), .z_share0(d0_P0_8_s0), .z_share1(d0_P0_8_s1));
  xor_module u_xor_P0_9_d0 (.x_share0(share0_in[9]), .x_share1(share1_in[9]), .y_share0(share0_in[41]), .y_share1(share1_in[41]), .z_share0(d0_P0_9_s0), .z_share1(d0_P0_9_s1));
  xor_module u_xor_o0_d0 (.x_share0(share0_in[0]), .x_share1(share1_in[0]), .y_share0(share0_in[32]), .y_share1(share1_in[32]), .z_share0(d0_o0_s0), .z_share1(d0_o0_s1));
  reg_module u_reg_P0_1_d1 (.clk(clk), .input_share0(d0_P0_1_s0), .input_share1(d0_P0_1_s1), .output_share0(d1_P0_1_s0), .output_share1(d1_P0_1_s1));
  reg_module u_reg_P0_10_d1 (.clk(clk), .input_share0(d0_P0_10_s0), .input_share1(d0_P0_10_s1), .output_share0(d1_P0_10_s0), .output_share1(d1_P0_10_s1));
  reg_module u_reg_P0_11_d1 (.clk(clk), .input_share0(d0_P0_11_s0), .input_share1(d0_P0_11_s1), .output_share0(d1_P0_11_s0), .output_share1(d1_P0_11_s1));
  reg_module u_reg_P0_12_d1 (.clk(clk), .input_share0(d0_P0_12_s0), .input_share1(d0_P0_12_s1), .output_share0(d1_P0_12_s0), .output_share1(d1_P0_12_s1));
  reg_module u_reg_P0_13_d1 (.clk(clk), .input_share0(d0_P0_13_s0), .input_share1(d0_P0_13_s1), .output_share0(d1_P0_13_s0), .output_share1(d1_P0_13_s1));
  reg_module u_reg_P0_14_d1 (.clk(clk), .input_share0(d0_P0_14_s0), .input_share1(d0_P0_14_s1), .output_share0(d1_P0_14_s0), .output_share1(d1_P0_14_s1));
  reg_module u_reg_P0_15_d1 (.clk(clk), .input_share0(d0_P0_15_s0), .input_share1(d0_P0_15_s1), .output_share0(d1_P0_15_s0), .output_share1(d1_P0_15_s1));
  reg_module u_reg_P0_16_d1 (.clk(clk), .input_share0(d0_P0_16_s0), .input_share1(d0_P0_16_s1), .output_share0(d1_P0_16_s0), .output_share1(d1_P0_16_s1));
  reg_module u_reg_P0_17_d1 (.clk(clk), .input_share0(d0_P0_17_s0), .input_share1(d0_P0_17_s1), .output_share0(d1_P0_17_s0), .output_share1(d1_P0_17_s1));
  reg_module u_reg_P0_18_d1 (.clk(clk), .input_share0(d0_P0_18_s0), .input_share1(d0_P0_18_s1), .output_share0(d1_P0_18_s0), .output_share1(d1_P0_18_s1));
  reg_module u_reg_P0_19_d1 (.clk(clk), .input_share0(d0_P0_19_s0), .input_share1(d0_P0_19_s1), .output_share0(d1_P0_19_s0), .output_share1(d1_P0_19_s1));
  reg_module u_reg_P0_2_d1 (.clk(clk), .input_share0(d0_P0_2_s0), .input_share1(d0_P0_2_s1), .output_share0(d1_P0_2_s0), .output_share1(d1_P0_2_s1));
  reg_module u_reg_P0_20_d1 (.clk(clk), .input_share0(d0_P0_20_s0), .input_share1(d0_P0_20_s1), .output_share0(d1_P0_20_s0), .output_share1(d1_P0_20_s1));
  reg_module u_reg_P0_21_d1 (.clk(clk), .input_share0(d0_P0_21_s0), .input_share1(d0_P0_21_s1), .output_share0(d1_P0_21_s0), .output_share1(d1_P0_21_s1));
  reg_module u_reg_P0_22_d1 (.clk(clk), .input_share0(d0_P0_22_s0), .input_share1(d0_P0_22_s1), .output_share0(d1_P0_22_s0), .output_share1(d1_P0_22_s1));
  reg_module u_reg_P0_23_d1 (.clk(clk), .input_share0(d0_P0_23_s0), .input_share1(d0_P0_23_s1), .output_share0(d1_P0_23_s0), .output_share1(d1_P0_23_s1));
  reg_module u_reg_P0_24_d1 (.clk(clk), .input_share0(d0_P0_24_s0), .input_share1(d0_P0_24_s1), .output_share0(d1_P0_24_s0), .output_share1(d1_P0_24_s1));
  reg_module u_reg_P0_25_d1 (.clk(clk), .input_share0(d0_P0_25_s0), .input_share1(d0_P0_25_s1), .output_share0(d1_P0_25_s0), .output_share1(d1_P0_25_s1));
  reg_module u_reg_P0_26_d1 (.clk(clk), .input_share0(d0_P0_26_s0), .input_share1(d0_P0_26_s1), .output_share0(d1_P0_26_s0), .output_share1(d1_P0_26_s1));
  reg_module u_reg_P0_27_d1 (.clk(clk), .input_share0(d0_P0_27_s0), .input_share1(d0_P0_27_s1), .output_share0(d1_P0_27_s0), .output_share1(d1_P0_27_s1));
  reg_module u_reg_P0_28_d1 (.clk(clk), .input_share0(d0_P0_28_s0), .input_share1(d0_P0_28_s1), .output_share0(d1_P0_28_s0), .output_share1(d1_P0_28_s1));
  reg_module u_reg_P0_29_d1 (.clk(clk), .input_share0(d0_P0_29_s0), .input_share1(d0_P0_29_s1), .output_share0(d1_P0_29_s0), .output_share1(d1_P0_29_s1));
  reg_module u_reg_P0_3_d1 (.clk(clk), .input_share0(d0_P0_3_s0), .input_share1(d0_P0_3_s1), .output_share0(d1_P0_3_s0), .output_share1(d1_P0_3_s1));
  reg_module u_reg_P0_30_d1 (.clk(clk), .input_share0(d0_P0_30_s0), .input_share1(d0_P0_30_s1), .output_share0(d1_P0_30_s0), .output_share1(d1_P0_30_s1));
  reg_module u_reg_P0_31_d1 (.clk(clk), .input_share0(d0_P0_31_s0), .input_share1(d0_P0_31_s1), .output_share0(d1_P0_31_s0), .output_share1(d1_P0_31_s1));
  reg_module u_reg_P0_4_d1 (.clk(clk), .input_share0(d0_P0_4_s0), .input_share1(d0_P0_4_s1), .output_share0(d1_P0_4_s0), .output_share1(d1_P0_4_s1));
  reg_module u_reg_P0_5_d1 (.clk(clk), .input_share0(d0_P0_5_s0), .input_share1(d0_P0_5_s1), .output_share0(d1_P0_5_s0), .output_share1(d1_P0_5_s1));
  reg_module u_reg_P0_6_d1 (.clk(clk), .input_share0(d0_P0_6_s0), .input_share1(d0_P0_6_s1), .output_share0(d1_P0_6_s0), .output_share1(d1_P0_6_s1));
  reg_module u_reg_P0_7_d1 (.clk(clk), .input_share0(d0_P0_7_s0), .input_share1(d0_P0_7_s1), .output_share0(d1_P0_7_s0), .output_share1(d1_P0_7_s1));
  reg_module u_reg_P0_8_d1 (.clk(clk), .input_share0(d0_P0_8_s0), .input_share1(d0_P0_8_s1), .output_share0(d1_P0_8_s0), .output_share1(d1_P0_8_s1));
  reg_module u_reg_P0_9_d1 (.clk(clk), .input_share0(d0_P0_9_s0), .input_share1(d0_P0_9_s1), .output_share0(d1_P0_9_s0), .output_share1(d1_P0_9_s1));
  and_module u_and_G0_0_d1 (.clk(clk), .x_share0(share0_in[0]), .x_share1(share1_in[0]), .y_share0(share0_in[32]), .y_share1(share1_in[32]), .rand(r_G0_0), .z_share0(d1_G0_0_s0), .z_share1(d1_G0_0_s1));
  assign r_G0_0 = rand_bit_share0[1];
  and_module u_and_G0_1_d1 (.clk(clk), .x_share0(share0_in[1]), .x_share1(share1_in[1]), .y_share0(share0_in[33]), .y_share1(share1_in[33]), .rand(r_G0_1), .z_share0(d1_G0_1_s0), .z_share1(d1_G0_1_s1));
  assign r_G0_1 = rand_bit_share0[0];
  and_module u_and_G0_10_d1 (.clk(clk), .x_share0(share0_in[10]), .x_share1(share1_in[10]), .y_share0(share0_in[42]), .y_share1(share1_in[42]), .rand(r_G0_10), .z_share0(d1_G0_10_s0), .z_share1(d1_G0_10_s1));
  assign r_G0_10 = rand_bit_share0[4];
  and_module u_and_G0_11_d1 (.clk(clk), .x_share0(share0_in[11]), .x_share1(share1_in[11]), .y_share0(share0_in[43]), .y_share1(share1_in[43]), .rand(r_G0_11), .z_share0(d1_G0_11_s0), .z_share1(d1_G0_11_s1));
  assign r_G0_11 = rand_bit_share0[2];
  and_module u_and_G0_12_d1 (.clk(clk), .x_share0(share0_in[12]), .x_share1(share1_in[12]), .y_share0(share0_in[44]), .y_share1(share1_in[44]), .rand(r_G0_12), .z_share0(d1_G0_12_s0), .z_share1(d1_G0_12_s1));
  assign r_G0_12 = rand_bit_share0[9];
  and_module u_and_G0_13_d1 (.clk(clk), .x_share0(share0_in[13]), .x_share1(share1_in[13]), .y_share0(share0_in[45]), .y_share1(share1_in[45]), .rand(r_G0_13), .z_share0(d1_G0_13_s0), .z_share1(d1_G0_13_s1));
  assign r_G0_13 = rand_bit_share0[0];
  and_module u_and_G0_14_d1 (.clk(clk), .x_share0(share0_in[14]), .x_share1(share1_in[14]), .y_share0(share0_in[46]), .y_share1(share1_in[46]), .rand(r_G0_14), .z_share0(d1_G0_14_s0), .z_share1(d1_G0_14_s1));
  assign r_G0_14 = rand_bit_share0[19];
  and_module u_and_G0_15_d1 (.clk(clk), .x_share0(share0_in[15]), .x_share1(share1_in[15]), .y_share0(share0_in[47]), .y_share1(share1_in[47]), .rand(r_G0_15), .z_share0(d1_G0_15_s0), .z_share1(d1_G0_15_s1));
  assign r_G0_15 = rand_bit_share0[1];
  and_module u_and_G0_16_d1 (.clk(clk), .x_share0(share0_in[16]), .x_share1(share1_in[16]), .y_share0(share0_in[48]), .y_share1(share1_in[48]), .rand(r_G0_16), .z_share0(d1_G0_16_s0), .z_share1(d1_G0_16_s1));
  assign r_G0_16 = rand_bit_share0[4];
  and_module u_and_G0_17_d1 (.clk(clk), .x_share0(share0_in[17]), .x_share1(share1_in[17]), .y_share0(share0_in[49]), .y_share1(share1_in[49]), .rand(r_G0_17), .z_share0(d1_G0_17_s0), .z_share1(d1_G0_17_s1));
  assign r_G0_17 = rand_bit_share0[2];
  and_module u_and_G0_18_d1 (.clk(clk), .x_share0(share0_in[18]), .x_share1(share1_in[18]), .y_share0(share0_in[50]), .y_share1(share1_in[50]), .rand(r_G0_18), .z_share0(d1_G0_18_s0), .z_share1(d1_G0_18_s1));
  assign r_G0_18 = rand_bit_share0[5];
  and_module u_and_G0_19_d1 (.clk(clk), .x_share0(share0_in[19]), .x_share1(share1_in[19]), .y_share0(share0_in[51]), .y_share1(share1_in[51]), .rand(r_G0_19), .z_share0(d1_G0_19_s0), .z_share1(d1_G0_19_s1));
  assign r_G0_19 = rand_bit_share0[0];
  and_module u_and_G0_2_d1 (.clk(clk), .x_share0(share0_in[2]), .x_share1(share1_in[2]), .y_share0(share0_in[34]), .y_share1(share1_in[34]), .rand(r_G0_2), .z_share0(d1_G0_2_s0), .z_share1(d1_G0_2_s1));
  assign r_G0_2 = rand_bit_share0[10];
  and_module u_and_G0_20_d1 (.clk(clk), .x_share0(share0_in[20]), .x_share1(share1_in[20]), .y_share0(share0_in[52]), .y_share1(share1_in[52]), .rand(r_G0_20), .z_share0(d1_G0_20_s0), .z_share1(d1_G0_20_s1));
  assign r_G0_20 = rand_bit_share0[3];
  and_module u_and_G0_21_d1 (.clk(clk), .x_share0(share0_in[21]), .x_share1(share1_in[21]), .y_share0(share0_in[53]), .y_share1(share1_in[53]), .rand(r_G0_21), .z_share0(d1_G0_21_s0), .z_share1(d1_G0_21_s1));
  assign r_G0_21 = rand_bit_share0[5];
  and_module u_and_G0_22_d1 (.clk(clk), .x_share0(share0_in[22]), .x_share1(share1_in[22]), .y_share0(share0_in[54]), .y_share1(share1_in[54]), .rand(r_G0_22), .z_share0(d1_G0_22_s0), .z_share1(d1_G0_22_s1));
  assign r_G0_22 = rand_bit_share0[1];
  and_module u_and_G0_23_d1 (.clk(clk), .x_share0(share0_in[23]), .x_share1(share1_in[23]), .y_share0(share0_in[55]), .y_share1(share1_in[55]), .rand(r_G0_23), .z_share0(d1_G0_23_s0), .z_share1(d1_G0_23_s1));
  assign r_G0_23 = rand_bit_share0[3];
  and_module u_and_G0_24_d1 (.clk(clk), .x_share0(share0_in[24]), .x_share1(share1_in[24]), .y_share0(share0_in[56]), .y_share1(share1_in[56]), .rand(r_G0_24), .z_share0(d1_G0_24_s0), .z_share1(d1_G0_24_s1));
  assign r_G0_24 = rand_bit_share0[2];
  and_module u_and_G0_25_d1 (.clk(clk), .x_share0(share0_in[25]), .x_share1(share1_in[25]), .y_share0(share0_in[57]), .y_share1(share1_in[57]), .rand(r_G0_25), .z_share0(d1_G0_25_s0), .z_share1(d1_G0_25_s1));
  assign r_G0_25 = rand_bit_share0[0];
  and_module u_and_G0_26_d1 (.clk(clk), .x_share0(share0_in[26]), .x_share1(share1_in[26]), .y_share0(share0_in[58]), .y_share1(share1_in[58]), .rand(r_G0_26), .z_share0(d1_G0_26_s0), .z_share1(d1_G0_26_s1));
  assign r_G0_26 = rand_bit_share0[9];
  and_module u_and_G0_27_d1 (.clk(clk), .x_share0(share0_in[27]), .x_share1(share1_in[27]), .y_share0(share0_in[59]), .y_share1(share1_in[59]), .rand(r_G0_27), .z_share0(d1_G0_27_s0), .z_share1(d1_G0_27_s1));
  assign r_G0_27 = rand_bit_share0[1];
  and_module u_and_G0_28_d1 (.clk(clk), .x_share0(share0_in[28]), .x_share1(share1_in[28]), .y_share0(share0_in[60]), .y_share1(share1_in[60]), .rand(r_G0_28), .z_share0(d1_G0_28_s0), .z_share1(d1_G0_28_s1));
  assign r_G0_28 = rand_bit_share0[4];
  and_module u_and_G0_29_d1 (.clk(clk), .x_share0(share0_in[29]), .x_share1(share1_in[29]), .y_share0(share0_in[61]), .y_share1(share1_in[61]), .rand(r_G0_29), .z_share0(d1_G0_29_s0), .z_share1(d1_G0_29_s1));
  assign r_G0_29 = rand_bit_share0[2];
  and_module u_and_G0_3_d1 (.clk(clk), .x_share0(share0_in[3]), .x_share1(share1_in[3]), .y_share0(share0_in[35]), .y_share1(share1_in[35]), .rand(r_G0_3), .z_share0(d1_G0_3_s0), .z_share1(d1_G0_3_s1));
  assign r_G0_3 = rand_bit_share0[1];
  and_module u_and_G0_30_d1 (.clk(clk), .x_share0(share0_in[30]), .x_share1(share1_in[30]), .y_share0(share0_in[62]), .y_share1(share1_in[62]), .rand(r_G0_30), .z_share0(d1_G0_30_s0), .z_share1(d1_G0_30_s1));
  assign r_G0_30 = rand_bit_share0[3];
  and_module u_and_G0_31_d1 (.clk(clk), .x_share0(share0_in[31]), .x_share1(share1_in[31]), .y_share0(share0_in[63]), .y_share1(share1_in[63]), .rand(r_G0_31), .z_share0(d1_G0_31_s0), .z_share1(d1_G0_31_s1));
  assign r_G0_31 = rand_bit_share0[0];
  and_module u_and_G0_4_d1 (.clk(clk), .x_share0(share0_in[4]), .x_share1(share1_in[4]), .y_share0(share0_in[36]), .y_share1(share1_in[36]), .rand(r_G0_4), .z_share0(d1_G0_4_s0), .z_share1(d1_G0_4_s1));
  assign r_G0_4 = rand_bit_share0[4];
  and_module u_and_G0_5_d1 (.clk(clk), .x_share0(share0_in[5]), .x_share1(share1_in[5]), .y_share0(share0_in[37]), .y_share1(share1_in[37]), .rand(r_G0_5), .z_share0(d1_G0_5_s0), .z_share1(d1_G0_5_s1));
  assign r_G0_5 = rand_bit_share0[2];
  and_module u_and_G0_6_d1 (.clk(clk), .x_share0(share0_in[6]), .x_share1(share1_in[6]), .y_share0(share0_in[38]), .y_share1(share1_in[38]), .rand(r_G0_6), .z_share0(d1_G0_6_s0), .z_share1(d1_G0_6_s1));
  assign r_G0_6 = rand_bit_share0[5];
  and_module u_and_G0_7_d1 (.clk(clk), .x_share0(share0_in[7]), .x_share1(share1_in[7]), .y_share0(share0_in[39]), .y_share1(share1_in[39]), .rand(r_G0_7), .z_share0(d1_G0_7_s0), .z_share1(d1_G0_7_s1));
  assign r_G0_7 = rand_bit_share0[0];
  and_module u_and_G0_8_d1 (.clk(clk), .x_share0(share0_in[8]), .x_share1(share1_in[8]), .y_share0(share0_in[40]), .y_share1(share1_in[40]), .rand(r_G0_8), .z_share0(d1_G0_8_s0), .z_share1(d1_G0_8_s1));
  assign r_G0_8 = rand_bit_share0[11];
  and_module u_and_G0_9_d1 (.clk(clk), .x_share0(share0_in[9]), .x_share1(share1_in[9]), .y_share0(share0_in[41]), .y_share1(share1_in[41]), .rand(r_G0_9), .z_share0(d1_G0_9_s0), .z_share1(d1_G0_9_s1));
  assign r_G0_9 = rand_bit_share0[1];
  and_module u_and_P1_10_d1 (.clk(clk), .x_share0(d0_P0_10_s0), .x_share1(d0_P0_10_s1), .y_share0(d0_P0_9_s0), .y_share1(d0_P0_9_s1), .rand(r_P1_10), .z_share0(d1_P1_10_s0), .z_share1(d1_P1_10_s1));
  assign r_P1_10 = rand_bit_share0[1];
  and_module u_and_P1_11_d1 (.clk(clk), .x_share0(d0_P0_11_s0), .x_share1(d0_P0_11_s1), .y_share0(d0_P0_10_s0), .y_share1(d0_P0_10_s1), .rand(r_P1_11), .z_share0(d1_P1_11_s0), .z_share1(d1_P1_11_s1));
  assign r_P1_11 = rand_bit_share0[7];
  and_module u_and_P1_12_d1 (.clk(clk), .x_share0(d0_P0_12_s0), .x_share1(d0_P0_12_s1), .y_share0(d0_P0_11_s0), .y_share1(d0_P0_11_s1), .rand(r_P1_12), .z_share0(d1_P1_12_s0), .z_share1(d1_P1_12_s1));
  assign r_P1_12 = rand_bit_share0[2];
  and_module u_and_P1_13_d1 (.clk(clk), .x_share0(d0_P0_13_s0), .x_share1(d0_P0_13_s1), .y_share0(d0_P0_12_s0), .y_share1(d0_P0_12_s1), .rand(r_P1_13), .z_share0(d1_P1_13_s0), .z_share1(d1_P1_13_s1));
  assign r_P1_13 = rand_bit_share0[6];
  and_module u_and_P1_14_d1 (.clk(clk), .x_share0(d0_P0_14_s0), .x_share1(d0_P0_14_s1), .y_share0(d0_P0_13_s0), .y_share1(d0_P0_13_s1), .rand(r_P1_14), .z_share0(d1_P1_14_s0), .z_share1(d1_P1_14_s1));
  assign r_P1_14 = rand_bit_share0[0];
  and_module u_and_P1_15_d1 (.clk(clk), .x_share0(d0_P0_15_s0), .x_share1(d0_P0_15_s1), .y_share0(d0_P0_14_s0), .y_share1(d0_P0_14_s1), .rand(r_P1_15), .z_share0(d1_P1_15_s0), .z_share1(d1_P1_15_s1));
  assign r_P1_15 = rand_bit_share0[8];
  and_module u_and_P1_16_d1 (.clk(clk), .x_share0(d0_P0_16_s0), .x_share1(d0_P0_16_s1), .y_share0(d0_P0_15_s0), .y_share1(d0_P0_15_s1), .rand(r_P1_16), .z_share0(d1_P1_16_s0), .z_share1(d1_P1_16_s1));
  assign r_P1_16 = rand_bit_share0[5];
  and_module u_and_P1_17_d1 (.clk(clk), .x_share0(d0_P0_17_s0), .x_share1(d0_P0_17_s1), .y_share0(d0_P0_16_s0), .y_share1(d0_P0_16_s1), .rand(r_P1_17), .z_share0(d1_P1_17_s0), .z_share1(d1_P1_17_s1));
  assign r_P1_17 = rand_bit_share0[3];
  and_module u_and_P1_18_d1 (.clk(clk), .x_share0(d0_P0_18_s0), .x_share1(d0_P0_18_s1), .y_share0(d0_P0_17_s0), .y_share1(d0_P0_17_s1), .rand(r_P1_18), .z_share0(d1_P1_18_s0), .z_share1(d1_P1_18_s1));
  assign r_P1_18 = rand_bit_share0[3];
  and_module u_and_P1_19_d1 (.clk(clk), .x_share0(d0_P0_19_s0), .x_share1(d0_P0_19_s1), .y_share0(d0_P0_18_s0), .y_share1(d0_P0_18_s1), .rand(r_P1_19), .z_share0(d1_P1_19_s0), .z_share1(d1_P1_19_s1));
  assign r_P1_19 = rand_bit_share0[5];
  and_module u_and_P1_2_d1 (.clk(clk), .x_share0(d0_P0_2_s0), .x_share1(d0_P0_2_s1), .y_share0(d0_P0_1_s0), .y_share1(d0_P0_1_s1), .rand(r_P1_2), .z_share0(d1_P1_2_s0), .z_share1(d1_P1_2_s1));
  assign r_P1_2 = rand_bit_share0[2];
  and_module u_and_P1_20_d1 (.clk(clk), .x_share0(d0_P0_20_s0), .x_share1(d0_P0_20_s1), .y_share0(d0_P0_19_s0), .y_share1(d0_P0_19_s1), .rand(r_P1_20), .z_share0(d1_P1_20_s0), .z_share1(d1_P1_20_s1));
  assign r_P1_20 = rand_bit_share0[1];
  and_module u_and_P1_21_d1 (.clk(clk), .x_share0(d0_P0_21_s0), .x_share1(d0_P0_21_s1), .y_share0(d0_P0_20_s0), .y_share1(d0_P0_20_s1), .rand(r_P1_21), .z_share0(d1_P1_21_s0), .z_share1(d1_P1_21_s1));
  assign r_P1_21 = rand_bit_share0[7];
  and_module u_and_P1_22_d1 (.clk(clk), .x_share0(d0_P0_22_s0), .x_share1(d0_P0_22_s1), .y_share0(d0_P0_21_s0), .y_share1(d0_P0_21_s1), .rand(r_P1_22), .z_share0(d1_P1_22_s0), .z_share1(d1_P1_22_s1));
  assign r_P1_22 = rand_bit_share0[2];
  and_module u_and_P1_23_d1 (.clk(clk), .x_share0(d0_P0_23_s0), .x_share1(d0_P0_23_s1), .y_share0(d0_P0_22_s0), .y_share1(d0_P0_22_s1), .rand(r_P1_23), .z_share0(d1_P1_23_s0), .z_share1(d1_P1_23_s1));
  assign r_P1_23 = rand_bit_share0[6];
  and_module u_and_P1_24_d1 (.clk(clk), .x_share0(d0_P0_24_s0), .x_share1(d0_P0_24_s1), .y_share0(d0_P0_23_s0), .y_share1(d0_P0_23_s1), .rand(r_P1_24), .z_share0(d1_P1_24_s0), .z_share1(d1_P1_24_s1));
  assign r_P1_24 = rand_bit_share0[0];
  and_module u_and_P1_25_d1 (.clk(clk), .x_share0(d0_P0_25_s0), .x_share1(d0_P0_25_s1), .y_share0(d0_P0_24_s0), .y_share1(d0_P0_24_s1), .rand(r_P1_25), .z_share0(d1_P1_25_s0), .z_share1(d1_P1_25_s1));
  assign r_P1_25 = rand_bit_share0[8];
  and_module u_and_P1_26_d1 (.clk(clk), .x_share0(d0_P0_26_s0), .x_share1(d0_P0_26_s1), .y_share0(d0_P0_25_s0), .y_share1(d0_P0_25_s1), .rand(r_P1_26), .z_share0(d1_P1_26_s0), .z_share1(d1_P1_26_s1));
  assign r_P1_26 = rand_bit_share0[12];
  and_module u_and_P1_27_d1 (.clk(clk), .x_share0(d0_P0_27_s0), .x_share1(d0_P0_27_s1), .y_share0(d0_P0_26_s0), .y_share1(d0_P0_26_s1), .rand(r_P1_27), .z_share0(d1_P1_27_s0), .z_share1(d1_P1_27_s1));
  assign r_P1_27 = rand_bit_share0[9];
  and_module u_and_P1_28_d1 (.clk(clk), .x_share0(d0_P0_28_s0), .x_share1(d0_P0_28_s1), .y_share0(d0_P0_27_s0), .y_share1(d0_P0_27_s1), .rand(r_P1_28), .z_share0(d1_P1_28_s0), .z_share1(d1_P1_28_s1));
  assign r_P1_28 = rand_bit_share0[8];
  and_module u_and_P1_29_d1 (.clk(clk), .x_share0(d0_P0_29_s0), .x_share1(d0_P0_29_s1), .y_share0(d0_P0_28_s0), .y_share1(d0_P0_28_s1), .rand(r_P1_29), .z_share0(d1_P1_29_s0), .z_share1(d1_P1_29_s1));
  assign r_P1_29 = rand_bit_share0[4];
  and_module u_and_P1_3_d1 (.clk(clk), .x_share0(d0_P0_3_s0), .x_share1(d0_P0_3_s1), .y_share0(d0_P0_2_s0), .y_share1(d0_P0_2_s1), .rand(r_P1_3), .z_share0(d1_P1_3_s0), .z_share1(d1_P1_3_s1));
  assign r_P1_3 = rand_bit_share0[15];
  and_module u_and_P1_30_d1 (.clk(clk), .x_share0(d0_P0_30_s0), .x_share1(d0_P0_30_s1), .y_share0(d0_P0_29_s0), .y_share1(d0_P0_29_s1), .rand(r_P1_30), .z_share0(d1_P1_30_s0), .z_share1(d1_P1_30_s1));
  assign r_P1_30 = rand_bit_share0[17];
  and_module u_and_P1_31_d1 (.clk(clk), .x_share0(d0_P0_31_s0), .x_share1(d0_P0_31_s1), .y_share0(d0_P0_30_s0), .y_share1(d0_P0_30_s1), .rand(r_P1_31), .z_share0(d1_P1_31_s0), .z_share1(d1_P1_31_s1));
  assign r_P1_31 = rand_bit_share0[14];
  and_module u_and_P1_4_d1 (.clk(clk), .x_share0(d0_P0_4_s0), .x_share1(d0_P0_4_s1), .y_share0(d0_P0_3_s0), .y_share1(d0_P0_3_s1), .rand(r_P1_4), .z_share0(d1_P1_4_s0), .z_share1(d1_P1_4_s1));
  assign r_P1_4 = rand_bit_share0[7];
  and_module u_and_P1_5_d1 (.clk(clk), .x_share0(d0_P0_5_s0), .x_share1(d0_P0_5_s1), .y_share0(d0_P0_4_s0), .y_share1(d0_P0_4_s1), .rand(r_P1_5), .z_share0(d1_P1_5_s0), .z_share1(d1_P1_5_s1));
  assign r_P1_5 = rand_bit_share0[14];
  and_module u_and_P1_6_d1 (.clk(clk), .x_share0(d0_P0_6_s0), .x_share1(d0_P0_6_s1), .y_share0(d0_P0_5_s0), .y_share1(d0_P0_5_s1), .rand(r_P1_6), .z_share0(d1_P1_6_s0), .z_share1(d1_P1_6_s1));
  assign r_P1_6 = rand_bit_share0[11];
  and_module u_and_P1_7_d1 (.clk(clk), .x_share0(d0_P0_7_s0), .x_share1(d0_P0_7_s1), .y_share0(d0_P0_6_s0), .y_share1(d0_P0_6_s1), .rand(r_P1_7), .z_share0(d1_P1_7_s0), .z_share1(d1_P1_7_s1));
  assign r_P1_7 = rand_bit_share0[12];
  and_module u_and_P1_8_d1 (.clk(clk), .x_share0(d0_P0_8_s0), .x_share1(d0_P0_8_s1), .y_share0(d0_P0_7_s0), .y_share1(d0_P0_7_s1), .rand(r_P1_8), .z_share0(d1_P1_8_s0), .z_share1(d1_P1_8_s1));
  assign r_P1_8 = rand_bit_share0[3];
  and_module u_and_P1_9_d1 (.clk(clk), .x_share0(d0_P0_9_s0), .x_share1(d0_P0_9_s1), .y_share0(d0_P0_8_s0), .y_share1(d0_P0_8_s1), .rand(r_P1_9), .z_share0(d1_P1_9_s0), .z_share1(d1_P1_9_s1));
  assign r_P1_9 = rand_bit_share0[9];
  xor_module u_xor_o1_d1 (.x_share0(d1_P0_1_s0), .x_share1(d1_P0_1_s1), .y_share0(d1_G0_0_s0), .y_share1(d1_G0_0_s1), .z_share0(d1_o1_s0), .z_share1(d1_o1_s1));
  reg_module u_reg_G0_0_d2 (.clk(clk), .input_share0(d1_G0_0_s0), .input_share1(d1_G0_0_s1), .output_share0(d2_G0_0_s0), .output_share1(d2_G0_0_s1));
  reg_module u_reg_G0_1_d2 (.clk(clk), .input_share0(d1_G0_1_s0), .input_share1(d1_G0_1_s1), .output_share0(d2_G0_1_s0), .output_share1(d2_G0_1_s1));
  reg_module u_reg_G0_10_d2 (.clk(clk), .input_share0(d1_G0_10_s0), .input_share1(d1_G0_10_s1), .output_share0(d2_G0_10_s0), .output_share1(d2_G0_10_s1));
  reg_module u_reg_G0_11_d2 (.clk(clk), .input_share0(d1_G0_11_s0), .input_share1(d1_G0_11_s1), .output_share0(d2_G0_11_s0), .output_share1(d2_G0_11_s1));
  reg_module u_reg_G0_12_d2 (.clk(clk), .input_share0(d1_G0_12_s0), .input_share1(d1_G0_12_s1), .output_share0(d2_G0_12_s0), .output_share1(d2_G0_12_s1));
  reg_module u_reg_G0_13_d2 (.clk(clk), .input_share0(d1_G0_13_s0), .input_share1(d1_G0_13_s1), .output_share0(d2_G0_13_s0), .output_share1(d2_G0_13_s1));
  reg_module u_reg_G0_14_d2 (.clk(clk), .input_share0(d1_G0_14_s0), .input_share1(d1_G0_14_s1), .output_share0(d2_G0_14_s0), .output_share1(d2_G0_14_s1));
  reg_module u_reg_G0_15_d2 (.clk(clk), .input_share0(d1_G0_15_s0), .input_share1(d1_G0_15_s1), .output_share0(d2_G0_15_s0), .output_share1(d2_G0_15_s1));
  reg_module u_reg_G0_16_d2 (.clk(clk), .input_share0(d1_G0_16_s0), .input_share1(d1_G0_16_s1), .output_share0(d2_G0_16_s0), .output_share1(d2_G0_16_s1));
  reg_module u_reg_G0_17_d2 (.clk(clk), .input_share0(d1_G0_17_s0), .input_share1(d1_G0_17_s1), .output_share0(d2_G0_17_s0), .output_share1(d2_G0_17_s1));
  reg_module u_reg_G0_18_d2 (.clk(clk), .input_share0(d1_G0_18_s0), .input_share1(d1_G0_18_s1), .output_share0(d2_G0_18_s0), .output_share1(d2_G0_18_s1));
  reg_module u_reg_G0_19_d2 (.clk(clk), .input_share0(d1_G0_19_s0), .input_share1(d1_G0_19_s1), .output_share0(d2_G0_19_s0), .output_share1(d2_G0_19_s1));
  reg_module u_reg_G0_2_d2 (.clk(clk), .input_share0(d1_G0_2_s0), .input_share1(d1_G0_2_s1), .output_share0(d2_G0_2_s0), .output_share1(d2_G0_2_s1));
  reg_module u_reg_G0_20_d2 (.clk(clk), .input_share0(d1_G0_20_s0), .input_share1(d1_G0_20_s1), .output_share0(d2_G0_20_s0), .output_share1(d2_G0_20_s1));
  reg_module u_reg_G0_21_d2 (.clk(clk), .input_share0(d1_G0_21_s0), .input_share1(d1_G0_21_s1), .output_share0(d2_G0_21_s0), .output_share1(d2_G0_21_s1));
  reg_module u_reg_G0_22_d2 (.clk(clk), .input_share0(d1_G0_22_s0), .input_share1(d1_G0_22_s1), .output_share0(d2_G0_22_s0), .output_share1(d2_G0_22_s1));
  reg_module u_reg_G0_23_d2 (.clk(clk), .input_share0(d1_G0_23_s0), .input_share1(d1_G0_23_s1), .output_share0(d2_G0_23_s0), .output_share1(d2_G0_23_s1));
  reg_module u_reg_G0_24_d2 (.clk(clk), .input_share0(d1_G0_24_s0), .input_share1(d1_G0_24_s1), .output_share0(d2_G0_24_s0), .output_share1(d2_G0_24_s1));
  reg_module u_reg_G0_25_d2 (.clk(clk), .input_share0(d1_G0_25_s0), .input_share1(d1_G0_25_s1), .output_share0(d2_G0_25_s0), .output_share1(d2_G0_25_s1));
  reg_module u_reg_G0_26_d2 (.clk(clk), .input_share0(d1_G0_26_s0), .input_share1(d1_G0_26_s1), .output_share0(d2_G0_26_s0), .output_share1(d2_G0_26_s1));
  reg_module u_reg_G0_27_d2 (.clk(clk), .input_share0(d1_G0_27_s0), .input_share1(d1_G0_27_s1), .output_share0(d2_G0_27_s0), .output_share1(d2_G0_27_s1));
  reg_module u_reg_G0_28_d2 (.clk(clk), .input_share0(d1_G0_28_s0), .input_share1(d1_G0_28_s1), .output_share0(d2_G0_28_s0), .output_share1(d2_G0_28_s1));
  reg_module u_reg_G0_29_d2 (.clk(clk), .input_share0(d1_G0_29_s0), .input_share1(d1_G0_29_s1), .output_share0(d2_G0_29_s0), .output_share1(d2_G0_29_s1));
  reg_module u_reg_G0_3_d2 (.clk(clk), .input_share0(d1_G0_3_s0), .input_share1(d1_G0_3_s1), .output_share0(d2_G0_3_s0), .output_share1(d2_G0_3_s1));
  reg_module u_reg_G0_30_d2 (.clk(clk), .input_share0(d1_G0_30_s0), .input_share1(d1_G0_30_s1), .output_share0(d2_G0_30_s0), .output_share1(d2_G0_30_s1));
  reg_module u_reg_G0_31_d2 (.clk(clk), .input_share0(d1_G0_31_s0), .input_share1(d1_G0_31_s1), .output_share0(d2_G0_31_s0), .output_share1(d2_G0_31_s1));
  reg_module u_reg_G0_4_d2 (.clk(clk), .input_share0(d1_G0_4_s0), .input_share1(d1_G0_4_s1), .output_share0(d2_G0_4_s0), .output_share1(d2_G0_4_s1));
  reg_module u_reg_G0_5_d2 (.clk(clk), .input_share0(d1_G0_5_s0), .input_share1(d1_G0_5_s1), .output_share0(d2_G0_5_s0), .output_share1(d2_G0_5_s1));
  reg_module u_reg_G0_6_d2 (.clk(clk), .input_share0(d1_G0_6_s0), .input_share1(d1_G0_6_s1), .output_share0(d2_G0_6_s0), .output_share1(d2_G0_6_s1));
  reg_module u_reg_G0_7_d2 (.clk(clk), .input_share0(d1_G0_7_s0), .input_share1(d1_G0_7_s1), .output_share0(d2_G0_7_s0), .output_share1(d2_G0_7_s1));
  reg_module u_reg_G0_8_d2 (.clk(clk), .input_share0(d1_G0_8_s0), .input_share1(d1_G0_8_s1), .output_share0(d2_G0_8_s0), .output_share1(d2_G0_8_s1));
  reg_module u_reg_G0_9_d2 (.clk(clk), .input_share0(d1_G0_9_s0), .input_share1(d1_G0_9_s1), .output_share0(d2_G0_9_s0), .output_share1(d2_G0_9_s1));
  reg_module u_reg_P0_10_d2 (.clk(clk), .input_share0(d1_P0_10_s0), .input_share1(d1_P0_10_s1), .output_share0(d2_P0_10_s0), .output_share1(d2_P0_10_s1));
  reg_module u_reg_P0_11_d2 (.clk(clk), .input_share0(d1_P0_11_s0), .input_share1(d1_P0_11_s1), .output_share0(d2_P0_11_s0), .output_share1(d2_P0_11_s1));
  reg_module u_reg_P0_12_d2 (.clk(clk), .input_share0(d1_P0_12_s0), .input_share1(d1_P0_12_s1), .output_share0(d2_P0_12_s0), .output_share1(d2_P0_12_s1));
  reg_module u_reg_P0_13_d2 (.clk(clk), .input_share0(d1_P0_13_s0), .input_share1(d1_P0_13_s1), .output_share0(d2_P0_13_s0), .output_share1(d2_P0_13_s1));
  reg_module u_reg_P0_14_d2 (.clk(clk), .input_share0(d1_P0_14_s0), .input_share1(d1_P0_14_s1), .output_share0(d2_P0_14_s0), .output_share1(d2_P0_14_s1));
  reg_module u_reg_P0_15_d2 (.clk(clk), .input_share0(d1_P0_15_s0), .input_share1(d1_P0_15_s1), .output_share0(d2_P0_15_s0), .output_share1(d2_P0_15_s1));
  reg_module u_reg_P0_16_d2 (.clk(clk), .input_share0(d1_P0_16_s0), .input_share1(d1_P0_16_s1), .output_share0(d2_P0_16_s0), .output_share1(d2_P0_16_s1));
  reg_module u_reg_P0_17_d2 (.clk(clk), .input_share0(d1_P0_17_s0), .input_share1(d1_P0_17_s1), .output_share0(d2_P0_17_s0), .output_share1(d2_P0_17_s1));
  reg_module u_reg_P0_18_d2 (.clk(clk), .input_share0(d1_P0_18_s0), .input_share1(d1_P0_18_s1), .output_share0(d2_P0_18_s0), .output_share1(d2_P0_18_s1));
  reg_module u_reg_P0_19_d2 (.clk(clk), .input_share0(d1_P0_19_s0), .input_share1(d1_P0_19_s1), .output_share0(d2_P0_19_s0), .output_share1(d2_P0_19_s1));
  reg_module u_reg_P0_2_d2 (.clk(clk), .input_share0(d1_P0_2_s0), .input_share1(d1_P0_2_s1), .output_share0(d2_P0_2_s0), .output_share1(d2_P0_2_s1));
  reg_module u_reg_P0_20_d2 (.clk(clk), .input_share0(d1_P0_20_s0), .input_share1(d1_P0_20_s1), .output_share0(d2_P0_20_s0), .output_share1(d2_P0_20_s1));
  reg_module u_reg_P0_21_d2 (.clk(clk), .input_share0(d1_P0_21_s0), .input_share1(d1_P0_21_s1), .output_share0(d2_P0_21_s0), .output_share1(d2_P0_21_s1));
  reg_module u_reg_P0_22_d2 (.clk(clk), .input_share0(d1_P0_22_s0), .input_share1(d1_P0_22_s1), .output_share0(d2_P0_22_s0), .output_share1(d2_P0_22_s1));
  reg_module u_reg_P0_23_d2 (.clk(clk), .input_share0(d1_P0_23_s0), .input_share1(d1_P0_23_s1), .output_share0(d2_P0_23_s0), .output_share1(d2_P0_23_s1));
  reg_module u_reg_P0_24_d2 (.clk(clk), .input_share0(d1_P0_24_s0), .input_share1(d1_P0_24_s1), .output_share0(d2_P0_24_s0), .output_share1(d2_P0_24_s1));
  reg_module u_reg_P0_25_d2 (.clk(clk), .input_share0(d1_P0_25_s0), .input_share1(d1_P0_25_s1), .output_share0(d2_P0_25_s0), .output_share1(d2_P0_25_s1));
  reg_module u_reg_P0_26_d2 (.clk(clk), .input_share0(d1_P0_26_s0), .input_share1(d1_P0_26_s1), .output_share0(d2_P0_26_s0), .output_share1(d2_P0_26_s1));
  reg_module u_reg_P0_27_d2 (.clk(clk), .input_share0(d1_P0_27_s0), .input_share1(d1_P0_27_s1), .output_share0(d2_P0_27_s0), .output_share1(d2_P0_27_s1));
  reg_module u_reg_P0_28_d2 (.clk(clk), .input_share0(d1_P0_28_s0), .input_share1(d1_P0_28_s1), .output_share0(d2_P0_28_s0), .output_share1(d2_P0_28_s1));
  reg_module u_reg_P0_29_d2 (.clk(clk), .input_share0(d1_P0_29_s0), .input_share1(d1_P0_29_s1), .output_share0(d2_P0_29_s0), .output_share1(d2_P0_29_s1));
  reg_module u_reg_P0_3_d2 (.clk(clk), .input_share0(d1_P0_3_s0), .input_share1(d1_P0_3_s1), .output_share0(d2_P0_3_s0), .output_share1(d2_P0_3_s1));
  reg_module u_reg_P0_30_d2 (.clk(clk), .input_share0(d1_P0_30_s0), .input_share1(d1_P0_30_s1), .output_share0(d2_P0_30_s0), .output_share1(d2_P0_30_s1));
  reg_module u_reg_P0_31_d2 (.clk(clk), .input_share0(d1_P0_31_s0), .input_share1(d1_P0_31_s1), .output_share0(d2_P0_31_s0), .output_share1(d2_P0_31_s1));
  reg_module u_reg_P0_4_d2 (.clk(clk), .input_share0(d1_P0_4_s0), .input_share1(d1_P0_4_s1), .output_share0(d2_P0_4_s0), .output_share1(d2_P0_4_s1));
  reg_module u_reg_P0_5_d2 (.clk(clk), .input_share0(d1_P0_5_s0), .input_share1(d1_P0_5_s1), .output_share0(d2_P0_5_s0), .output_share1(d2_P0_5_s1));
  reg_module u_reg_P0_6_d2 (.clk(clk), .input_share0(d1_P0_6_s0), .input_share1(d1_P0_6_s1), .output_share0(d2_P0_6_s0), .output_share1(d2_P0_6_s1));
  reg_module u_reg_P0_7_d2 (.clk(clk), .input_share0(d1_P0_7_s0), .input_share1(d1_P0_7_s1), .output_share0(d2_P0_7_s0), .output_share1(d2_P0_7_s1));
  reg_module u_reg_P0_8_d2 (.clk(clk), .input_share0(d1_P0_8_s0), .input_share1(d1_P0_8_s1), .output_share0(d2_P0_8_s0), .output_share1(d2_P0_8_s1));
  reg_module u_reg_P0_9_d2 (.clk(clk), .input_share0(d1_P0_9_s0), .input_share1(d1_P0_9_s1), .output_share0(d2_P0_9_s0), .output_share1(d2_P0_9_s1));
  reg_module u_reg_P1_10_d2 (.clk(clk), .input_share0(d1_P1_10_s0), .input_share1(d1_P1_10_s1), .output_share0(d2_P1_10_s0), .output_share1(d2_P1_10_s1));
  reg_module u_reg_P1_11_d2 (.clk(clk), .input_share0(d1_P1_11_s0), .input_share1(d1_P1_11_s1), .output_share0(d2_P1_11_s0), .output_share1(d2_P1_11_s1));
  reg_module u_reg_P1_12_d2 (.clk(clk), .input_share0(d1_P1_12_s0), .input_share1(d1_P1_12_s1), .output_share0(d2_P1_12_s0), .output_share1(d2_P1_12_s1));
  reg_module u_reg_P1_13_d2 (.clk(clk), .input_share0(d1_P1_13_s0), .input_share1(d1_P1_13_s1), .output_share0(d2_P1_13_s0), .output_share1(d2_P1_13_s1));
  reg_module u_reg_P1_14_d2 (.clk(clk), .input_share0(d1_P1_14_s0), .input_share1(d1_P1_14_s1), .output_share0(d2_P1_14_s0), .output_share1(d2_P1_14_s1));
  reg_module u_reg_P1_15_d2 (.clk(clk), .input_share0(d1_P1_15_s0), .input_share1(d1_P1_15_s1), .output_share0(d2_P1_15_s0), .output_share1(d2_P1_15_s1));
  reg_module u_reg_P1_16_d2 (.clk(clk), .input_share0(d1_P1_16_s0), .input_share1(d1_P1_16_s1), .output_share0(d2_P1_16_s0), .output_share1(d2_P1_16_s1));
  reg_module u_reg_P1_17_d2 (.clk(clk), .input_share0(d1_P1_17_s0), .input_share1(d1_P1_17_s1), .output_share0(d2_P1_17_s0), .output_share1(d2_P1_17_s1));
  reg_module u_reg_P1_18_d2 (.clk(clk), .input_share0(d1_P1_18_s0), .input_share1(d1_P1_18_s1), .output_share0(d2_P1_18_s0), .output_share1(d2_P1_18_s1));
  reg_module u_reg_P1_19_d2 (.clk(clk), .input_share0(d1_P1_19_s0), .input_share1(d1_P1_19_s1), .output_share0(d2_P1_19_s0), .output_share1(d2_P1_19_s1));
  reg_module u_reg_P1_20_d2 (.clk(clk), .input_share0(d1_P1_20_s0), .input_share1(d1_P1_20_s1), .output_share0(d2_P1_20_s0), .output_share1(d2_P1_20_s1));
  reg_module u_reg_P1_21_d2 (.clk(clk), .input_share0(d1_P1_21_s0), .input_share1(d1_P1_21_s1), .output_share0(d2_P1_21_s0), .output_share1(d2_P1_21_s1));
  reg_module u_reg_P1_22_d2 (.clk(clk), .input_share0(d1_P1_22_s0), .input_share1(d1_P1_22_s1), .output_share0(d2_P1_22_s0), .output_share1(d2_P1_22_s1));
  reg_module u_reg_P1_23_d2 (.clk(clk), .input_share0(d1_P1_23_s0), .input_share1(d1_P1_23_s1), .output_share0(d2_P1_23_s0), .output_share1(d2_P1_23_s1));
  reg_module u_reg_P1_24_d2 (.clk(clk), .input_share0(d1_P1_24_s0), .input_share1(d1_P1_24_s1), .output_share0(d2_P1_24_s0), .output_share1(d2_P1_24_s1));
  reg_module u_reg_P1_25_d2 (.clk(clk), .input_share0(d1_P1_25_s0), .input_share1(d1_P1_25_s1), .output_share0(d2_P1_25_s0), .output_share1(d2_P1_25_s1));
  reg_module u_reg_P1_26_d2 (.clk(clk), .input_share0(d1_P1_26_s0), .input_share1(d1_P1_26_s1), .output_share0(d2_P1_26_s0), .output_share1(d2_P1_26_s1));
  reg_module u_reg_P1_27_d2 (.clk(clk), .input_share0(d1_P1_27_s0), .input_share1(d1_P1_27_s1), .output_share0(d2_P1_27_s0), .output_share1(d2_P1_27_s1));
  reg_module u_reg_P1_28_d2 (.clk(clk), .input_share0(d1_P1_28_s0), .input_share1(d1_P1_28_s1), .output_share0(d2_P1_28_s0), .output_share1(d2_P1_28_s1));
  reg_module u_reg_P1_29_d2 (.clk(clk), .input_share0(d1_P1_29_s0), .input_share1(d1_P1_29_s1), .output_share0(d2_P1_29_s0), .output_share1(d2_P1_29_s1));
  reg_module u_reg_P1_3_d2 (.clk(clk), .input_share0(d1_P1_3_s0), .input_share1(d1_P1_3_s1), .output_share0(d2_P1_3_s0), .output_share1(d2_P1_3_s1));
  reg_module u_reg_P1_30_d2 (.clk(clk), .input_share0(d1_P1_30_s0), .input_share1(d1_P1_30_s1), .output_share0(d2_P1_30_s0), .output_share1(d2_P1_30_s1));
  reg_module u_reg_P1_31_d2 (.clk(clk), .input_share0(d1_P1_31_s0), .input_share1(d1_P1_31_s1), .output_share0(d2_P1_31_s0), .output_share1(d2_P1_31_s1));
  reg_module u_reg_P1_4_d2 (.clk(clk), .input_share0(d1_P1_4_s0), .input_share1(d1_P1_4_s1), .output_share0(d2_P1_4_s0), .output_share1(d2_P1_4_s1));
  reg_module u_reg_P1_5_d2 (.clk(clk), .input_share0(d1_P1_5_s0), .input_share1(d1_P1_5_s1), .output_share0(d2_P1_5_s0), .output_share1(d2_P1_5_s1));
  reg_module u_reg_P1_6_d2 (.clk(clk), .input_share0(d1_P1_6_s0), .input_share1(d1_P1_6_s1), .output_share0(d2_P1_6_s0), .output_share1(d2_P1_6_s1));
  reg_module u_reg_P1_7_d2 (.clk(clk), .input_share0(d1_P1_7_s0), .input_share1(d1_P1_7_s1), .output_share0(d2_P1_7_s0), .output_share1(d2_P1_7_s1));
  reg_module u_reg_P1_8_d2 (.clk(clk), .input_share0(d1_P1_8_s0), .input_share1(d1_P1_8_s1), .output_share0(d2_P1_8_s0), .output_share1(d2_P1_8_s1));
  reg_module u_reg_P1_9_d2 (.clk(clk), .input_share0(d1_P1_9_s0), .input_share1(d1_P1_9_s1), .output_share0(d2_P1_9_s0), .output_share1(d2_P1_9_s1));
  xor_module u_xor_G1_1_d2 (.x_share0(d2_t0_s0), .x_share1(d2_t0_s1), .y_share0(d2_G0_1_s0), .y_share1(d2_G0_1_s1), .z_share0(d2_G1_1_s0), .z_share1(d2_G1_1_s1));
  xor_module u_xor_G1_10_d2 (.x_share0(d2_t9_s0), .x_share1(d2_t9_s1), .y_share0(d2_G0_10_s0), .y_share1(d2_G0_10_s1), .z_share0(d2_G1_10_s0), .z_share1(d2_G1_10_s1));
  xor_module u_xor_G1_11_d2 (.x_share0(d2_t10_s0), .x_share1(d2_t10_s1), .y_share0(d2_G0_11_s0), .y_share1(d2_G0_11_s1), .z_share0(d2_G1_11_s0), .z_share1(d2_G1_11_s1));
  xor_module u_xor_G1_12_d2 (.x_share0(d2_t11_s0), .x_share1(d2_t11_s1), .y_share0(d2_G0_12_s0), .y_share1(d2_G0_12_s1), .z_share0(d2_G1_12_s0), .z_share1(d2_G1_12_s1));
  xor_module u_xor_G1_13_d2 (.x_share0(d2_t12_s0), .x_share1(d2_t12_s1), .y_share0(d2_G0_13_s0), .y_share1(d2_G0_13_s1), .z_share0(d2_G1_13_s0), .z_share1(d2_G1_13_s1));
  xor_module u_xor_G1_14_d2 (.x_share0(d2_t13_s0), .x_share1(d2_t13_s1), .y_share0(d2_G0_14_s0), .y_share1(d2_G0_14_s1), .z_share0(d2_G1_14_s0), .z_share1(d2_G1_14_s1));
  xor_module u_xor_G1_15_d2 (.x_share0(d2_t14_s0), .x_share1(d2_t14_s1), .y_share0(d2_G0_15_s0), .y_share1(d2_G0_15_s1), .z_share0(d2_G1_15_s0), .z_share1(d2_G1_15_s1));
  xor_module u_xor_G1_16_d2 (.x_share0(d2_t15_s0), .x_share1(d2_t15_s1), .y_share0(d2_G0_16_s0), .y_share1(d2_G0_16_s1), .z_share0(d2_G1_16_s0), .z_share1(d2_G1_16_s1));
  xor_module u_xor_G1_17_d2 (.x_share0(d2_t16_s0), .x_share1(d2_t16_s1), .y_share0(d2_G0_17_s0), .y_share1(d2_G0_17_s1), .z_share0(d2_G1_17_s0), .z_share1(d2_G1_17_s1));
  xor_module u_xor_G1_18_d2 (.x_share0(d2_t17_s0), .x_share1(d2_t17_s1), .y_share0(d2_G0_18_s0), .y_share1(d2_G0_18_s1), .z_share0(d2_G1_18_s0), .z_share1(d2_G1_18_s1));
  xor_module u_xor_G1_19_d2 (.x_share0(d2_t18_s0), .x_share1(d2_t18_s1), .y_share0(d2_G0_19_s0), .y_share1(d2_G0_19_s1), .z_share0(d2_G1_19_s0), .z_share1(d2_G1_19_s1));
  xor_module u_xor_G1_2_d2 (.x_share0(d2_t1_s0), .x_share1(d2_t1_s1), .y_share0(d2_G0_2_s0), .y_share1(d2_G0_2_s1), .z_share0(d2_G1_2_s0), .z_share1(d2_G1_2_s1));
  xor_module u_xor_G1_20_d2 (.x_share0(d2_t19_s0), .x_share1(d2_t19_s1), .y_share0(d2_G0_20_s0), .y_share1(d2_G0_20_s1), .z_share0(d2_G1_20_s0), .z_share1(d2_G1_20_s1));
  xor_module u_xor_G1_21_d2 (.x_share0(d2_t20_s0), .x_share1(d2_t20_s1), .y_share0(d2_G0_21_s0), .y_share1(d2_G0_21_s1), .z_share0(d2_G1_21_s0), .z_share1(d2_G1_21_s1));
  xor_module u_xor_G1_22_d2 (.x_share0(d2_t21_s0), .x_share1(d2_t21_s1), .y_share0(d2_G0_22_s0), .y_share1(d2_G0_22_s1), .z_share0(d2_G1_22_s0), .z_share1(d2_G1_22_s1));
  xor_module u_xor_G1_23_d2 (.x_share0(d2_t22_s0), .x_share1(d2_t22_s1), .y_share0(d2_G0_23_s0), .y_share1(d2_G0_23_s1), .z_share0(d2_G1_23_s0), .z_share1(d2_G1_23_s1));
  xor_module u_xor_G1_24_d2 (.x_share0(d2_t23_s0), .x_share1(d2_t23_s1), .y_share0(d2_G0_24_s0), .y_share1(d2_G0_24_s1), .z_share0(d2_G1_24_s0), .z_share1(d2_G1_24_s1));
  xor_module u_xor_G1_25_d2 (.x_share0(d2_t24_s0), .x_share1(d2_t24_s1), .y_share0(d2_G0_25_s0), .y_share1(d2_G0_25_s1), .z_share0(d2_G1_25_s0), .z_share1(d2_G1_25_s1));
  xor_module u_xor_G1_26_d2 (.x_share0(d2_t25_s0), .x_share1(d2_t25_s1), .y_share0(d2_G0_26_s0), .y_share1(d2_G0_26_s1), .z_share0(d2_G1_26_s0), .z_share1(d2_G1_26_s1));
  xor_module u_xor_G1_27_d2 (.x_share0(d2_t26_s0), .x_share1(d2_t26_s1), .y_share0(d2_G0_27_s0), .y_share1(d2_G0_27_s1), .z_share0(d2_G1_27_s0), .z_share1(d2_G1_27_s1));
  xor_module u_xor_G1_28_d2 (.x_share0(d2_t27_s0), .x_share1(d2_t27_s1), .y_share0(d2_G0_28_s0), .y_share1(d2_G0_28_s1), .z_share0(d2_G1_28_s0), .z_share1(d2_G1_28_s1));
  xor_module u_xor_G1_29_d2 (.x_share0(d2_t28_s0), .x_share1(d2_t28_s1), .y_share0(d2_G0_29_s0), .y_share1(d2_G0_29_s1), .z_share0(d2_G1_29_s0), .z_share1(d2_G1_29_s1));
  xor_module u_xor_G1_3_d2 (.x_share0(d2_t2_s0), .x_share1(d2_t2_s1), .y_share0(d2_G0_3_s0), .y_share1(d2_G0_3_s1), .z_share0(d2_G1_3_s0), .z_share1(d2_G1_3_s1));
  xor_module u_xor_G1_30_d2 (.x_share0(d2_t29_s0), .x_share1(d2_t29_s1), .y_share0(d2_G0_30_s0), .y_share1(d2_G0_30_s1), .z_share0(d2_G1_30_s0), .z_share1(d2_G1_30_s1));
  xor_module u_xor_G1_31_d2 (.x_share0(d2_t30_s0), .x_share1(d2_t30_s1), .y_share0(d2_G0_31_s0), .y_share1(d2_G0_31_s1), .z_share0(d2_G1_31_s0), .z_share1(d2_G1_31_s1));
  xor_module u_xor_G1_4_d2 (.x_share0(d2_t3_s0), .x_share1(d2_t3_s1), .y_share0(d2_G0_4_s0), .y_share1(d2_G0_4_s1), .z_share0(d2_G1_4_s0), .z_share1(d2_G1_4_s1));
  xor_module u_xor_G1_5_d2 (.x_share0(d2_t4_s0), .x_share1(d2_t4_s1), .y_share0(d2_G0_5_s0), .y_share1(d2_G0_5_s1), .z_share0(d2_G1_5_s0), .z_share1(d2_G1_5_s1));
  xor_module u_xor_G1_6_d2 (.x_share0(d2_t5_s0), .x_share1(d2_t5_s1), .y_share0(d2_G0_6_s0), .y_share1(d2_G0_6_s1), .z_share0(d2_G1_6_s0), .z_share1(d2_G1_6_s1));
  xor_module u_xor_G1_7_d2 (.x_share0(d2_t6_s0), .x_share1(d2_t6_s1), .y_share0(d2_G0_7_s0), .y_share1(d2_G0_7_s1), .z_share0(d2_G1_7_s0), .z_share1(d2_G1_7_s1));
  xor_module u_xor_G1_8_d2 (.x_share0(d2_t7_s0), .x_share1(d2_t7_s1), .y_share0(d2_G0_8_s0), .y_share1(d2_G0_8_s1), .z_share0(d2_G1_8_s0), .z_share1(d2_G1_8_s1));
  xor_module u_xor_G1_9_d2 (.x_share0(d2_t8_s0), .x_share1(d2_t8_s1), .y_share0(d2_G0_9_s0), .y_share1(d2_G0_9_s1), .z_share0(d2_G1_9_s0), .z_share1(d2_G1_9_s1));
  xor_module u_xor_G2_2_d2 (.x_share0(d2_t31_s0), .x_share1(d2_t31_s1), .y_share0(d2_G1_2_s0), .y_share1(d2_G1_2_s1), .z_share0(d2_G2_2_s0), .z_share1(d2_G2_2_s1));
  and_module u_and_P2_10_d2 (.clk(clk), .x_share0(d1_P1_10_s0), .x_share1(d1_P1_10_s1), .y_share0(d1_P1_8_s0), .y_share1(d1_P1_8_s1), .rand(r_P2_10), .z_share0(d2_P2_10_s0), .z_share1(d2_P2_10_s1));
  assign r_P2_10 = stage2_share0[17];
  and_module u_and_P2_11_d2 (.clk(clk), .x_share0(d1_P1_11_s0), .x_share1(d1_P1_11_s1), .y_share0(d1_P1_9_s0), .y_share1(d1_P1_9_s1), .rand(r_P2_11), .z_share0(d2_P2_11_s0), .z_share1(d2_P2_11_s1));
  assign r_P2_11 = stage2_share0[20];
  and_module u_and_P2_12_d2 (.clk(clk), .x_share0(d1_P1_12_s0), .x_share1(d1_P1_12_s1), .y_share0(d1_P1_10_s0), .y_share1(d1_P1_10_s1), .rand(r_P2_12), .z_share0(d2_P2_12_s0), .z_share1(d2_P2_12_s1));
  assign r_P2_12 = stage2_share0[14];
  and_module u_and_P2_13_d2 (.clk(clk), .x_share0(d1_P1_13_s0), .x_share1(d1_P1_13_s1), .y_share0(d1_P1_11_s0), .y_share1(d1_P1_11_s1), .rand(r_P2_13), .z_share0(d2_P2_13_s0), .z_share1(d2_P2_13_s1));
  assign r_P2_13 = stage2_share0[15];
  and_module u_and_P2_14_d2 (.clk(clk), .x_share0(d1_P1_14_s0), .x_share1(d1_P1_14_s1), .y_share0(d1_P1_12_s0), .y_share1(d1_P1_12_s1), .rand(r_P2_14), .z_share0(d2_P2_14_s0), .z_share1(d2_P2_14_s1));
  assign r_P2_14 = stage2_share0[7];
  and_module u_and_P2_15_d2 (.clk(clk), .x_share0(d1_P1_15_s0), .x_share1(d1_P1_15_s1), .y_share0(d1_P1_13_s0), .y_share1(d1_P1_13_s1), .rand(r_P2_15), .z_share0(d2_P2_15_s0), .z_share1(d2_P2_15_s1));
  assign r_P2_15 = stage2_share0[18];
  and_module u_and_P2_16_d2 (.clk(clk), .x_share0(d1_P1_16_s0), .x_share1(d1_P1_16_s1), .y_share0(d1_P1_14_s0), .y_share1(d1_P1_14_s1), .rand(r_P2_16), .z_share0(d2_P2_16_s0), .z_share1(d2_P2_16_s1));
  assign r_P2_16 = stage2_share0[23];
  and_module u_and_P2_17_d2 (.clk(clk), .x_share0(d1_P1_17_s0), .x_share1(d1_P1_17_s1), .y_share0(d1_P1_15_s0), .y_share1(d1_P1_15_s1), .rand(r_P2_17), .z_share0(d2_P2_17_s0), .z_share1(d2_P2_17_s1));
  assign r_P2_17 = stage2_share0[16];
  and_module u_and_P2_18_d2 (.clk(clk), .x_share0(d1_P1_18_s0), .x_share1(d1_P1_18_s1), .y_share0(d1_P1_16_s0), .y_share1(d1_P1_16_s1), .rand(r_P2_18), .z_share0(d2_P2_18_s0), .z_share1(d2_P2_18_s1));
  assign r_P2_18 = stage2_share0[8];
  and_module u_and_P2_19_d2 (.clk(clk), .x_share0(d1_P1_19_s0), .x_share1(d1_P1_19_s1), .y_share0(d1_P1_17_s0), .y_share1(d1_P1_17_s1), .rand(r_P2_19), .z_share0(d2_P2_19_s0), .z_share1(d2_P2_19_s1));
  assign r_P2_19 = stage2_share0[13];
  and_module u_and_P2_20_d2 (.clk(clk), .x_share0(d1_P1_20_s0), .x_share1(d1_P1_20_s1), .y_share0(d1_P1_18_s0), .y_share1(d1_P1_18_s1), .rand(r_P2_20), .z_share0(d2_P2_20_s0), .z_share1(d2_P2_20_s1));
  assign r_P2_20 = stage2_share0[13];
  and_module u_and_P2_21_d2 (.clk(clk), .x_share0(d1_P1_21_s0), .x_share1(d1_P1_21_s1), .y_share0(d1_P1_19_s0), .y_share1(d1_P1_19_s1), .rand(r_P2_21), .z_share0(d2_P2_21_s0), .z_share1(d2_P2_21_s1));
  assign r_P2_21 = stage2_share0[17];
  and_module u_and_P2_22_d2 (.clk(clk), .x_share0(d1_P1_22_s0), .x_share1(d1_P1_22_s1), .y_share0(d1_P1_20_s0), .y_share1(d1_P1_20_s1), .rand(r_P2_22), .z_share0(d2_P2_22_s0), .z_share1(d2_P2_22_s1));
  assign r_P2_22 = stage2_share0[10];
  and_module u_and_P2_23_d2 (.clk(clk), .x_share0(d1_P1_23_s0), .x_share1(d1_P1_23_s1), .y_share0(d1_P1_21_s0), .y_share1(d1_P1_21_s1), .rand(r_P2_23), .z_share0(d2_P2_23_s0), .z_share1(d2_P2_23_s1));
  assign r_P2_23 = stage2_share0[11];
  and_module u_and_P2_24_d2 (.clk(clk), .x_share0(d1_P1_24_s0), .x_share1(d1_P1_24_s1), .y_share0(d1_P1_22_s0), .y_share1(d1_P1_22_s1), .rand(r_P2_24), .z_share0(d2_P2_24_s0), .z_share1(d2_P2_24_s1));
  assign r_P2_24 = stage2_share0[18];
  and_module u_and_P2_25_d2 (.clk(clk), .x_share0(d1_P1_25_s0), .x_share1(d1_P1_25_s1), .y_share0(d1_P1_23_s0), .y_share1(d1_P1_23_s1), .rand(r_P2_25), .z_share0(d2_P2_25_s0), .z_share1(d2_P2_25_s1));
  assign r_P2_25 = stage2_share0[18];
  and_module u_and_P2_26_d2 (.clk(clk), .x_share0(d1_P1_26_s0), .x_share1(d1_P1_26_s1), .y_share0(d1_P1_24_s0), .y_share1(d1_P1_24_s1), .rand(r_P2_26), .z_share0(d2_P2_26_s0), .z_share1(d2_P2_26_s1));
  assign r_P2_26 = stage2_share0[15];
  and_module u_and_P2_27_d2 (.clk(clk), .x_share0(d1_P1_27_s0), .x_share1(d1_P1_27_s1), .y_share0(d1_P1_25_s0), .y_share1(d1_P1_25_s1), .rand(r_P2_27), .z_share0(d2_P2_27_s0), .z_share1(d2_P2_27_s1));
  assign r_P2_27 = stage2_share0[10];
  and_module u_and_P2_28_d2 (.clk(clk), .x_share0(d1_P1_28_s0), .x_share1(d1_P1_28_s1), .y_share0(d1_P1_26_s0), .y_share1(d1_P1_26_s1), .rand(r_P2_28), .z_share0(d2_P2_28_s0), .z_share1(d2_P2_28_s1));
  assign r_P2_28 = stage2_share0[19];
  and_module u_and_P2_29_d2 (.clk(clk), .x_share0(d1_P1_29_s0), .x_share1(d1_P1_29_s1), .y_share0(d1_P1_27_s0), .y_share1(d1_P1_27_s1), .rand(r_P2_29), .z_share0(d2_P2_29_s0), .z_share1(d2_P2_29_s1));
  assign r_P2_29 = stage2_share0[21];
  and_module u_and_P2_30_d2 (.clk(clk), .x_share0(d1_P1_30_s0), .x_share1(d1_P1_30_s1), .y_share0(d1_P1_28_s0), .y_share1(d1_P1_28_s1), .rand(r_P2_30), .z_share0(d2_P2_30_s0), .z_share1(d2_P2_30_s1));
  assign r_P2_30 = stage2_share0[18];
  and_module u_and_P2_31_d2 (.clk(clk), .x_share0(d1_P1_31_s0), .x_share1(d1_P1_31_s1), .y_share0(d1_P1_29_s0), .y_share1(d1_P1_29_s1), .rand(r_P2_31), .z_share0(d2_P2_31_s0), .z_share1(d2_P2_31_s1));
  assign r_P2_31 = stage2_share0[20];
  and_module u_and_P2_4_d2 (.clk(clk), .x_share0(d1_P1_4_s0), .x_share1(d1_P1_4_s1), .y_share0(d1_P1_2_s0), .y_share1(d1_P1_2_s1), .rand(r_P2_4), .z_share0(d2_P2_4_s0), .z_share1(d2_P2_4_s1));
  assign r_P2_4 = stage2_share0[0];
  and_module u_and_P2_5_d2 (.clk(clk), .x_share0(d1_P1_5_s0), .x_share1(d1_P1_5_s1), .y_share0(d1_P1_3_s0), .y_share1(d1_P1_3_s1), .rand(r_P2_5), .z_share0(d2_P2_5_s0), .z_share1(d2_P2_5_s1));
  assign r_P2_5 = stage2_share0[8];
  and_module u_and_P2_6_d2 (.clk(clk), .x_share0(d1_P1_6_s0), .x_share1(d1_P1_6_s1), .y_share0(d1_P1_4_s0), .y_share1(d1_P1_4_s1), .rand(r_P2_6), .z_share0(d2_P2_6_s0), .z_share1(d2_P2_6_s1));
  assign r_P2_6 = stage2_share0[12];
  and_module u_and_P2_7_d2 (.clk(clk), .x_share0(d1_P1_7_s0), .x_share1(d1_P1_7_s1), .y_share0(d1_P1_5_s0), .y_share1(d1_P1_5_s1), .rand(r_P2_7), .z_share0(d2_P2_7_s0), .z_share1(d2_P2_7_s1));
  assign r_P2_7 = stage2_share0[2];
  and_module u_and_P2_8_d2 (.clk(clk), .x_share0(d1_P1_8_s0), .x_share1(d1_P1_8_s1), .y_share0(d1_P1_6_s0), .y_share1(d1_P1_6_s1), .rand(r_P2_8), .z_share0(d2_P2_8_s0), .z_share1(d2_P2_8_s1));
  assign r_P2_8 = stage2_share0[9];
  and_module u_and_P2_9_d2 (.clk(clk), .x_share0(d1_P1_9_s0), .x_share1(d1_P1_9_s1), .y_share0(d1_P1_7_s0), .y_share1(d1_P1_7_s1), .rand(r_P2_9), .z_share0(d2_P2_9_s0), .z_share1(d2_P2_9_s1));
  assign r_P2_9 = stage2_share0[11];
  xor_module u_xor_o2_d2 (.x_share0(d2_P0_2_s0), .x_share1(d2_P0_2_s1), .y_share0(d2_G1_1_s0), .y_share1(d2_G1_1_s1), .z_share0(d2_o2_s0), .z_share1(d2_o2_s1));
  xor_module u_xor_o3_d2 (.x_share0(d2_P0_3_s0), .x_share1(d2_P0_3_s1), .y_share0(d2_G2_2_s0), .y_share1(d2_G2_2_s1), .z_share0(d2_o3_s0), .z_share1(d2_o3_s1));
  and_module u_and_t0_d2 (.clk(clk), .x_share0(d1_P0_1_s0), .x_share1(d1_P0_1_s1), .y_share0(d1_G0_0_s0), .y_share1(d1_G0_0_s1), .rand(r_t0), .z_share0(d2_t0_s0), .z_share1(d2_t0_s1));
  assign r_t0 = stage2_share0[5];
  and_module u_and_t1_d2 (.clk(clk), .x_share0(d1_P0_2_s0), .x_share1(d1_P0_2_s1), .y_share0(d1_G0_1_s0), .y_share1(d1_G0_1_s1), .rand(r_t1), .z_share0(d2_t1_s0), .z_share1(d2_t1_s1));
  assign r_t1 = stage2_share0[20];
  and_module u_and_t10_d2 (.clk(clk), .x_share0(d1_P0_11_s0), .x_share1(d1_P0_11_s1), .y_share0(d1_G0_10_s0), .y_share1(d1_G0_10_s1), .rand(r_t10), .z_share0(d2_t10_s0), .z_share1(d2_t10_s1));
  assign r_t10 = stage2_share0[14];
  and_module u_and_t11_d2 (.clk(clk), .x_share0(d1_P0_12_s0), .x_share1(d1_P0_12_s1), .y_share0(d1_G0_11_s0), .y_share1(d1_G0_11_s1), .rand(r_t11), .z_share0(d2_t11_s0), .z_share1(d2_t11_s1));
  assign r_t11 = stage2_share0[10];
  and_module u_and_t12_d2 (.clk(clk), .x_share0(d1_P0_13_s0), .x_share1(d1_P0_13_s1), .y_share0(d1_G0_12_s0), .y_share1(d1_G0_12_s1), .rand(r_t12), .z_share0(d2_t12_s0), .z_share1(d2_t12_s1));
  assign r_t12 = stage2_share0[11];
  and_module u_and_t13_d2 (.clk(clk), .x_share0(d1_P0_14_s0), .x_share1(d1_P0_14_s1), .y_share0(d1_G0_13_s0), .y_share1(d1_G0_13_s1), .rand(r_t13), .z_share0(d2_t13_s0), .z_share1(d2_t13_s1));
  assign r_t13 = stage2_share0[20];
  and_module u_and_t14_d2 (.clk(clk), .x_share0(d1_P0_15_s0), .x_share1(d1_P0_15_s1), .y_share0(d1_G0_14_s0), .y_share1(d1_G0_14_s1), .rand(r_t14), .z_share0(d2_t14_s0), .z_share1(d2_t14_s1));
  assign r_t14 = stage2_share0[4];
  and_module u_and_t15_d2 (.clk(clk), .x_share0(d1_P0_16_s0), .x_share1(d1_P0_16_s1), .y_share0(d1_G0_15_s0), .y_share1(d1_G0_15_s1), .rand(r_t15), .z_share0(d2_t15_s0), .z_share1(d2_t15_s1));
  assign r_t15 = stage2_share0[6];
  and_module u_and_t16_d2 (.clk(clk), .x_share0(d1_P0_17_s0), .x_share1(d1_P0_17_s1), .y_share0(d1_G0_16_s0), .y_share1(d1_G0_16_s1), .rand(r_t16), .z_share0(d2_t16_s0), .z_share1(d2_t16_s1));
  assign r_t16 = stage2_share0[14];
  and_module u_and_t17_d2 (.clk(clk), .x_share0(d1_P0_18_s0), .x_share1(d1_P0_18_s1), .y_share0(d1_G0_17_s0), .y_share1(d1_G0_17_s1), .rand(r_t17), .z_share0(d2_t17_s0), .z_share1(d2_t17_s1));
  assign r_t17 = stage2_share0[11];
  and_module u_and_t18_d2 (.clk(clk), .x_share0(d1_P0_19_s0), .x_share1(d1_P0_19_s1), .y_share0(d1_G0_18_s0), .y_share1(d1_G0_18_s1), .rand(r_t18), .z_share0(d2_t18_s0), .z_share1(d2_t18_s1));
  assign r_t18 = stage2_share0[12];
  and_module u_and_t19_d2 (.clk(clk), .x_share0(d1_P0_20_s0), .x_share1(d1_P0_20_s1), .y_share0(d1_G0_19_s0), .y_share1(d1_G0_19_s1), .rand(r_t19), .z_share0(d2_t19_s0), .z_share1(d2_t19_s1));
  assign r_t19 = stage2_share0[16];
  and_module u_and_t2_d2 (.clk(clk), .x_share0(d1_P0_3_s0), .x_share1(d1_P0_3_s1), .y_share0(d1_G0_2_s0), .y_share1(d1_G0_2_s1), .rand(r_t2), .z_share0(d2_t2_s0), .z_share1(d2_t2_s1));
  assign r_t2 = stage2_share0[4];
  and_module u_and_t20_d2 (.clk(clk), .x_share0(d1_P0_21_s0), .x_share1(d1_P0_21_s1), .y_share0(d1_G0_20_s0), .y_share1(d1_G0_20_s1), .rand(r_t20), .z_share0(d2_t20_s0), .z_share1(d2_t20_s1));
  assign r_t20 = stage2_share0[1];
  and_module u_and_t21_d2 (.clk(clk), .x_share0(d1_P0_22_s0), .x_share1(d1_P0_22_s1), .y_share0(d1_G0_21_s0), .y_share1(d1_G0_21_s1), .rand(r_t21), .z_share0(d2_t21_s0), .z_share1(d2_t21_s1));
  assign r_t21 = stage2_share0[4];
  and_module u_and_t22_d2 (.clk(clk), .x_share0(d1_P0_23_s0), .x_share1(d1_P0_23_s1), .y_share0(d1_G0_22_s0), .y_share1(d1_G0_22_s1), .rand(r_t22), .z_share0(d2_t22_s0), .z_share1(d2_t22_s1));
  assign r_t22 = stage2_share0[7];
  and_module u_and_t23_d2 (.clk(clk), .x_share0(d1_P0_24_s0), .x_share1(d1_P0_24_s1), .y_share0(d1_G0_23_s0), .y_share1(d1_G0_23_s1), .rand(r_t23), .z_share0(d2_t23_s0), .z_share1(d2_t23_s1));
  assign r_t23 = stage2_share0[14];
  and_module u_and_t24_d2 (.clk(clk), .x_share0(d1_P0_25_s0), .x_share1(d1_P0_25_s1), .y_share0(d1_G0_24_s0), .y_share1(d1_G0_24_s1), .rand(r_t24), .z_share0(d2_t24_s0), .z_share1(d2_t24_s1));
  assign r_t24 = stage2_share0[6];
  and_module u_and_t25_d2 (.clk(clk), .x_share0(d1_P0_26_s0), .x_share1(d1_P0_26_s1), .y_share0(d1_G0_25_s0), .y_share1(d1_G0_25_s1), .rand(r_t25), .z_share0(d2_t25_s0), .z_share1(d2_t25_s1));
  assign r_t25 = stage2_share0[10];
  and_module u_and_t26_d2 (.clk(clk), .x_share0(d1_P0_27_s0), .x_share1(d1_P0_27_s1), .y_share0(d1_G0_26_s0), .y_share1(d1_G0_26_s1), .rand(r_t26), .z_share0(d2_t26_s0), .z_share1(d2_t26_s1));
  assign r_t26 = stage2_share0[15];
  and_module u_and_t27_d2 (.clk(clk), .x_share0(d1_P0_28_s0), .x_share1(d1_P0_28_s1), .y_share0(d1_G0_27_s0), .y_share1(d1_G0_27_s1), .rand(r_t27), .z_share0(d2_t27_s0), .z_share1(d2_t27_s1));
  assign r_t27 = stage2_share0[7];
  and_module u_and_t28_d2 (.clk(clk), .x_share0(d1_P0_29_s0), .x_share1(d1_P0_29_s1), .y_share0(d1_G0_28_s0), .y_share1(d1_G0_28_s1), .rand(r_t28), .z_share0(d2_t28_s0), .z_share1(d2_t28_s1));
  assign r_t28 = stage2_share0[12];
  and_module u_and_t29_d2 (.clk(clk), .x_share0(d1_P0_30_s0), .x_share1(d1_P0_30_s1), .y_share0(d1_G0_29_s0), .y_share1(d1_G0_29_s1), .rand(r_t29), .z_share0(d2_t29_s0), .z_share1(d2_t29_s1));
  assign r_t29 = stage2_share0[5];
  and_module u_and_t3_d2 (.clk(clk), .x_share0(d1_P0_4_s0), .x_share1(d1_P0_4_s1), .y_share0(d1_G0_3_s0), .y_share1(d1_G0_3_s1), .rand(r_t3), .z_share0(d2_t3_s0), .z_share1(d2_t3_s1));
  assign r_t3 = stage2_share0[6];
  and_module u_and_t30_d2 (.clk(clk), .x_share0(d1_P0_31_s0), .x_share1(d1_P0_31_s1), .y_share0(d1_G0_30_s0), .y_share1(d1_G0_30_s1), .rand(r_t30), .z_share0(d2_t30_s0), .z_share1(d2_t30_s1));
  assign r_t30 = stage2_share0[16];
  and_module u_and_t31_d2 (.clk(clk), .x_share0(d1_P1_2_s0), .x_share1(d1_P1_2_s1), .y_share0(d1_G0_0_s0), .y_share1(d1_G0_0_s1), .rand(r_t31), .z_share0(d2_t31_s0), .z_share1(d2_t31_s1));
  assign r_t31 = stage2_share0[21];
  and_module u_and_t4_d2 (.clk(clk), .x_share0(d1_P0_5_s0), .x_share1(d1_P0_5_s1), .y_share0(d1_G0_4_s0), .y_share1(d1_G0_4_s1), .rand(r_t4), .z_share0(d2_t4_s0), .z_share1(d2_t4_s1));
  assign r_t4 = stage2_share0[13];
  and_module u_and_t5_d2 (.clk(clk), .x_share0(d1_P0_6_s0), .x_share1(d1_P0_6_s1), .y_share0(d1_G0_5_s0), .y_share1(d1_G0_5_s1), .rand(r_t5), .z_share0(d2_t5_s0), .z_share1(d2_t5_s1));
  assign r_t5 = stage2_share0[13];
  and_module u_and_t6_d2 (.clk(clk), .x_share0(d1_P0_7_s0), .x_share1(d1_P0_7_s1), .y_share0(d1_G0_6_s0), .y_share1(d1_G0_6_s1), .rand(r_t6), .z_share0(d2_t6_s0), .z_share1(d2_t6_s1));
  assign r_t6 = stage2_share0[16];
  and_module u_and_t7_d2 (.clk(clk), .x_share0(d1_P0_8_s0), .x_share1(d1_P0_8_s1), .y_share0(d1_G0_7_s0), .y_share1(d1_G0_7_s1), .rand(r_t7), .z_share0(d2_t7_s0), .z_share1(d2_t7_s1));
  assign r_t7 = stage2_share0[12];
  and_module u_and_t8_d2 (.clk(clk), .x_share0(d1_P0_9_s0), .x_share1(d1_P0_9_s1), .y_share0(d1_G0_8_s0), .y_share1(d1_G0_8_s1), .rand(r_t8), .z_share0(d2_t8_s0), .z_share1(d2_t8_s1));
  assign r_t8 = stage2_share0[10];
  and_module u_and_t9_d2 (.clk(clk), .x_share0(d1_P0_10_s0), .x_share1(d1_P0_10_s1), .y_share0(d1_G0_9_s0), .y_share1(d1_G0_9_s1), .rand(r_t9), .z_share0(d2_t9_s0), .z_share1(d2_t9_s1));
  assign r_t9 = stage2_share0[6];
  reg_module u_reg_G0_0_d3 (.clk(clk), .input_share0(d2_G0_0_s0), .input_share1(d2_G0_0_s1), .output_share0(d3_G0_0_s0), .output_share1(d3_G0_0_s1));
  reg_module u_reg_G1_1_d3 (.clk(clk), .input_share0(d2_G1_1_s0), .input_share1(d2_G1_1_s1), .output_share0(d3_G1_1_s0), .output_share1(d3_G1_1_s1));
  reg_module u_reg_G1_10_d3 (.clk(clk), .input_share0(d2_G1_10_s0), .input_share1(d2_G1_10_s1), .output_share0(d3_G1_10_s0), .output_share1(d3_G1_10_s1));
  reg_module u_reg_G1_11_d3 (.clk(clk), .input_share0(d2_G1_11_s0), .input_share1(d2_G1_11_s1), .output_share0(d3_G1_11_s0), .output_share1(d3_G1_11_s1));
  reg_module u_reg_G1_12_d3 (.clk(clk), .input_share0(d2_G1_12_s0), .input_share1(d2_G1_12_s1), .output_share0(d3_G1_12_s0), .output_share1(d3_G1_12_s1));
  reg_module u_reg_G1_13_d3 (.clk(clk), .input_share0(d2_G1_13_s0), .input_share1(d2_G1_13_s1), .output_share0(d3_G1_13_s0), .output_share1(d3_G1_13_s1));
  reg_module u_reg_G1_14_d3 (.clk(clk), .input_share0(d2_G1_14_s0), .input_share1(d2_G1_14_s1), .output_share0(d3_G1_14_s0), .output_share1(d3_G1_14_s1));
  reg_module u_reg_G1_15_d3 (.clk(clk), .input_share0(d2_G1_15_s0), .input_share1(d2_G1_15_s1), .output_share0(d3_G1_15_s0), .output_share1(d3_G1_15_s1));
  reg_module u_reg_G1_16_d3 (.clk(clk), .input_share0(d2_G1_16_s0), .input_share1(d2_G1_16_s1), .output_share0(d3_G1_16_s0), .output_share1(d3_G1_16_s1));
  reg_module u_reg_G1_17_d3 (.clk(clk), .input_share0(d2_G1_17_s0), .input_share1(d2_G1_17_s1), .output_share0(d3_G1_17_s0), .output_share1(d3_G1_17_s1));
  reg_module u_reg_G1_18_d3 (.clk(clk), .input_share0(d2_G1_18_s0), .input_share1(d2_G1_18_s1), .output_share0(d3_G1_18_s0), .output_share1(d3_G1_18_s1));
  reg_module u_reg_G1_19_d3 (.clk(clk), .input_share0(d2_G1_19_s0), .input_share1(d2_G1_19_s1), .output_share0(d3_G1_19_s0), .output_share1(d3_G1_19_s1));
  reg_module u_reg_G1_20_d3 (.clk(clk), .input_share0(d2_G1_20_s0), .input_share1(d2_G1_20_s1), .output_share0(d3_G1_20_s0), .output_share1(d3_G1_20_s1));
  reg_module u_reg_G1_21_d3 (.clk(clk), .input_share0(d2_G1_21_s0), .input_share1(d2_G1_21_s1), .output_share0(d3_G1_21_s0), .output_share1(d3_G1_21_s1));
  reg_module u_reg_G1_22_d3 (.clk(clk), .input_share0(d2_G1_22_s0), .input_share1(d2_G1_22_s1), .output_share0(d3_G1_22_s0), .output_share1(d3_G1_22_s1));
  reg_module u_reg_G1_23_d3 (.clk(clk), .input_share0(d2_G1_23_s0), .input_share1(d2_G1_23_s1), .output_share0(d3_G1_23_s0), .output_share1(d3_G1_23_s1));
  reg_module u_reg_G1_24_d3 (.clk(clk), .input_share0(d2_G1_24_s0), .input_share1(d2_G1_24_s1), .output_share0(d3_G1_24_s0), .output_share1(d3_G1_24_s1));
  reg_module u_reg_G1_25_d3 (.clk(clk), .input_share0(d2_G1_25_s0), .input_share1(d2_G1_25_s1), .output_share0(d3_G1_25_s0), .output_share1(d3_G1_25_s1));
  reg_module u_reg_G1_26_d3 (.clk(clk), .input_share0(d2_G1_26_s0), .input_share1(d2_G1_26_s1), .output_share0(d3_G1_26_s0), .output_share1(d3_G1_26_s1));
  reg_module u_reg_G1_27_d3 (.clk(clk), .input_share0(d2_G1_27_s0), .input_share1(d2_G1_27_s1), .output_share0(d3_G1_27_s0), .output_share1(d3_G1_27_s1));
  reg_module u_reg_G1_28_d3 (.clk(clk), .input_share0(d2_G1_28_s0), .input_share1(d2_G1_28_s1), .output_share0(d3_G1_28_s0), .output_share1(d3_G1_28_s1));
  reg_module u_reg_G1_29_d3 (.clk(clk), .input_share0(d2_G1_29_s0), .input_share1(d2_G1_29_s1), .output_share0(d3_G1_29_s0), .output_share1(d3_G1_29_s1));
  reg_module u_reg_G1_3_d3 (.clk(clk), .input_share0(d2_G1_3_s0), .input_share1(d2_G1_3_s1), .output_share0(d3_G1_3_s0), .output_share1(d3_G1_3_s1));
  reg_module u_reg_G1_30_d3 (.clk(clk), .input_share0(d2_G1_30_s0), .input_share1(d2_G1_30_s1), .output_share0(d3_G1_30_s0), .output_share1(d3_G1_30_s1));
  reg_module u_reg_G1_31_d3 (.clk(clk), .input_share0(d2_G1_31_s0), .input_share1(d2_G1_31_s1), .output_share0(d3_G1_31_s0), .output_share1(d3_G1_31_s1));
  reg_module u_reg_G1_4_d3 (.clk(clk), .input_share0(d2_G1_4_s0), .input_share1(d2_G1_4_s1), .output_share0(d3_G1_4_s0), .output_share1(d3_G1_4_s1));
  reg_module u_reg_G1_5_d3 (.clk(clk), .input_share0(d2_G1_5_s0), .input_share1(d2_G1_5_s1), .output_share0(d3_G1_5_s0), .output_share1(d3_G1_5_s1));
  reg_module u_reg_G1_6_d3 (.clk(clk), .input_share0(d2_G1_6_s0), .input_share1(d2_G1_6_s1), .output_share0(d3_G1_6_s0), .output_share1(d3_G1_6_s1));
  reg_module u_reg_G1_7_d3 (.clk(clk), .input_share0(d2_G1_7_s0), .input_share1(d2_G1_7_s1), .output_share0(d3_G1_7_s0), .output_share1(d3_G1_7_s1));
  reg_module u_reg_G1_8_d3 (.clk(clk), .input_share0(d2_G1_8_s0), .input_share1(d2_G1_8_s1), .output_share0(d3_G1_8_s0), .output_share1(d3_G1_8_s1));
  reg_module u_reg_G1_9_d3 (.clk(clk), .input_share0(d2_G1_9_s0), .input_share1(d2_G1_9_s1), .output_share0(d3_G1_9_s0), .output_share1(d3_G1_9_s1));
  reg_module u_reg_G2_2_d3 (.clk(clk), .input_share0(d2_G2_2_s0), .input_share1(d2_G2_2_s1), .output_share0(d3_G2_2_s0), .output_share1(d3_G2_2_s1));
  reg_module u_reg_P0_10_d3 (.clk(clk), .input_share0(d2_P0_10_s0), .input_share1(d2_P0_10_s1), .output_share0(d3_P0_10_s0), .output_share1(d3_P0_10_s1));
  reg_module u_reg_P0_11_d3 (.clk(clk), .input_share0(d2_P0_11_s0), .input_share1(d2_P0_11_s1), .output_share0(d3_P0_11_s0), .output_share1(d3_P0_11_s1));
  reg_module u_reg_P0_12_d3 (.clk(clk), .input_share0(d2_P0_12_s0), .input_share1(d2_P0_12_s1), .output_share0(d3_P0_12_s0), .output_share1(d3_P0_12_s1));
  reg_module u_reg_P0_13_d3 (.clk(clk), .input_share0(d2_P0_13_s0), .input_share1(d2_P0_13_s1), .output_share0(d3_P0_13_s0), .output_share1(d3_P0_13_s1));
  reg_module u_reg_P0_14_d3 (.clk(clk), .input_share0(d2_P0_14_s0), .input_share1(d2_P0_14_s1), .output_share0(d3_P0_14_s0), .output_share1(d3_P0_14_s1));
  reg_module u_reg_P0_15_d3 (.clk(clk), .input_share0(d2_P0_15_s0), .input_share1(d2_P0_15_s1), .output_share0(d3_P0_15_s0), .output_share1(d3_P0_15_s1));
  reg_module u_reg_P0_16_d3 (.clk(clk), .input_share0(d2_P0_16_s0), .input_share1(d2_P0_16_s1), .output_share0(d3_P0_16_s0), .output_share1(d3_P0_16_s1));
  reg_module u_reg_P0_17_d3 (.clk(clk), .input_share0(d2_P0_17_s0), .input_share1(d2_P0_17_s1), .output_share0(d3_P0_17_s0), .output_share1(d3_P0_17_s1));
  reg_module u_reg_P0_18_d3 (.clk(clk), .input_share0(d2_P0_18_s0), .input_share1(d2_P0_18_s1), .output_share0(d3_P0_18_s0), .output_share1(d3_P0_18_s1));
  reg_module u_reg_P0_19_d3 (.clk(clk), .input_share0(d2_P0_19_s0), .input_share1(d2_P0_19_s1), .output_share0(d3_P0_19_s0), .output_share1(d3_P0_19_s1));
  reg_module u_reg_P0_20_d3 (.clk(clk), .input_share0(d2_P0_20_s0), .input_share1(d2_P0_20_s1), .output_share0(d3_P0_20_s0), .output_share1(d3_P0_20_s1));
  reg_module u_reg_P0_21_d3 (.clk(clk), .input_share0(d2_P0_21_s0), .input_share1(d2_P0_21_s1), .output_share0(d3_P0_21_s0), .output_share1(d3_P0_21_s1));
  reg_module u_reg_P0_22_d3 (.clk(clk), .input_share0(d2_P0_22_s0), .input_share1(d2_P0_22_s1), .output_share0(d3_P0_22_s0), .output_share1(d3_P0_22_s1));
  reg_module u_reg_P0_23_d3 (.clk(clk), .input_share0(d2_P0_23_s0), .input_share1(d2_P0_23_s1), .output_share0(d3_P0_23_s0), .output_share1(d3_P0_23_s1));
  reg_module u_reg_P0_24_d3 (.clk(clk), .input_share0(d2_P0_24_s0), .input_share1(d2_P0_24_s1), .output_share0(d3_P0_24_s0), .output_share1(d3_P0_24_s1));
  reg_module u_reg_P0_25_d3 (.clk(clk), .input_share0(d2_P0_25_s0), .input_share1(d2_P0_25_s1), .output_share0(d3_P0_25_s0), .output_share1(d3_P0_25_s1));
  reg_module u_reg_P0_26_d3 (.clk(clk), .input_share0(d2_P0_26_s0), .input_share1(d2_P0_26_s1), .output_share0(d3_P0_26_s0), .output_share1(d3_P0_26_s1));
  reg_module u_reg_P0_27_d3 (.clk(clk), .input_share0(d2_P0_27_s0), .input_share1(d2_P0_27_s1), .output_share0(d3_P0_27_s0), .output_share1(d3_P0_27_s1));
  reg_module u_reg_P0_28_d3 (.clk(clk), .input_share0(d2_P0_28_s0), .input_share1(d2_P0_28_s1), .output_share0(d3_P0_28_s0), .output_share1(d3_P0_28_s1));
  reg_module u_reg_P0_29_d3 (.clk(clk), .input_share0(d2_P0_29_s0), .input_share1(d2_P0_29_s1), .output_share0(d3_P0_29_s0), .output_share1(d3_P0_29_s1));
  reg_module u_reg_P0_30_d3 (.clk(clk), .input_share0(d2_P0_30_s0), .input_share1(d2_P0_30_s1), .output_share0(d3_P0_30_s0), .output_share1(d3_P0_30_s1));
  reg_module u_reg_P0_31_d3 (.clk(clk), .input_share0(d2_P0_31_s0), .input_share1(d2_P0_31_s1), .output_share0(d3_P0_31_s0), .output_share1(d3_P0_31_s1));
  reg_module u_reg_P0_4_d3 (.clk(clk), .input_share0(d2_P0_4_s0), .input_share1(d2_P0_4_s1), .output_share0(d3_P0_4_s0), .output_share1(d3_P0_4_s1));
  reg_module u_reg_P0_5_d3 (.clk(clk), .input_share0(d2_P0_5_s0), .input_share1(d2_P0_5_s1), .output_share0(d3_P0_5_s0), .output_share1(d3_P0_5_s1));
  reg_module u_reg_P0_6_d3 (.clk(clk), .input_share0(d2_P0_6_s0), .input_share1(d2_P0_6_s1), .output_share0(d3_P0_6_s0), .output_share1(d3_P0_6_s1));
  reg_module u_reg_P0_7_d3 (.clk(clk), .input_share0(d2_P0_7_s0), .input_share1(d2_P0_7_s1), .output_share0(d3_P0_7_s0), .output_share1(d3_P0_7_s1));
  reg_module u_reg_P0_8_d3 (.clk(clk), .input_share0(d2_P0_8_s0), .input_share1(d2_P0_8_s1), .output_share0(d3_P0_8_s0), .output_share1(d3_P0_8_s1));
  reg_module u_reg_P0_9_d3 (.clk(clk), .input_share0(d2_P0_9_s0), .input_share1(d2_P0_9_s1), .output_share0(d3_P0_9_s0), .output_share1(d3_P0_9_s1));
  reg_module u_reg_P2_10_d3 (.clk(clk), .input_share0(d2_P2_10_s0), .input_share1(d2_P2_10_s1), .output_share0(d3_P2_10_s0), .output_share1(d3_P2_10_s1));
  reg_module u_reg_P2_11_d3 (.clk(clk), .input_share0(d2_P2_11_s0), .input_share1(d2_P2_11_s1), .output_share0(d3_P2_11_s0), .output_share1(d3_P2_11_s1));
  reg_module u_reg_P2_12_d3 (.clk(clk), .input_share0(d2_P2_12_s0), .input_share1(d2_P2_12_s1), .output_share0(d3_P2_12_s0), .output_share1(d3_P2_12_s1));
  reg_module u_reg_P2_13_d3 (.clk(clk), .input_share0(d2_P2_13_s0), .input_share1(d2_P2_13_s1), .output_share0(d3_P2_13_s0), .output_share1(d3_P2_13_s1));
  reg_module u_reg_P2_14_d3 (.clk(clk), .input_share0(d2_P2_14_s0), .input_share1(d2_P2_14_s1), .output_share0(d3_P2_14_s0), .output_share1(d3_P2_14_s1));
  reg_module u_reg_P2_15_d3 (.clk(clk), .input_share0(d2_P2_15_s0), .input_share1(d2_P2_15_s1), .output_share0(d3_P2_15_s0), .output_share1(d3_P2_15_s1));
  reg_module u_reg_P2_16_d3 (.clk(clk), .input_share0(d2_P2_16_s0), .input_share1(d2_P2_16_s1), .output_share0(d3_P2_16_s0), .output_share1(d3_P2_16_s1));
  reg_module u_reg_P2_17_d3 (.clk(clk), .input_share0(d2_P2_17_s0), .input_share1(d2_P2_17_s1), .output_share0(d3_P2_17_s0), .output_share1(d3_P2_17_s1));
  reg_module u_reg_P2_18_d3 (.clk(clk), .input_share0(d2_P2_18_s0), .input_share1(d2_P2_18_s1), .output_share0(d3_P2_18_s0), .output_share1(d3_P2_18_s1));
  reg_module u_reg_P2_19_d3 (.clk(clk), .input_share0(d2_P2_19_s0), .input_share1(d2_P2_19_s1), .output_share0(d3_P2_19_s0), .output_share1(d3_P2_19_s1));
  reg_module u_reg_P2_20_d3 (.clk(clk), .input_share0(d2_P2_20_s0), .input_share1(d2_P2_20_s1), .output_share0(d3_P2_20_s0), .output_share1(d3_P2_20_s1));
  reg_module u_reg_P2_21_d3 (.clk(clk), .input_share0(d2_P2_21_s0), .input_share1(d2_P2_21_s1), .output_share0(d3_P2_21_s0), .output_share1(d3_P2_21_s1));
  reg_module u_reg_P2_22_d3 (.clk(clk), .input_share0(d2_P2_22_s0), .input_share1(d2_P2_22_s1), .output_share0(d3_P2_22_s0), .output_share1(d3_P2_22_s1));
  reg_module u_reg_P2_23_d3 (.clk(clk), .input_share0(d2_P2_23_s0), .input_share1(d2_P2_23_s1), .output_share0(d3_P2_23_s0), .output_share1(d3_P2_23_s1));
  reg_module u_reg_P2_24_d3 (.clk(clk), .input_share0(d2_P2_24_s0), .input_share1(d2_P2_24_s1), .output_share0(d3_P2_24_s0), .output_share1(d3_P2_24_s1));
  reg_module u_reg_P2_25_d3 (.clk(clk), .input_share0(d2_P2_25_s0), .input_share1(d2_P2_25_s1), .output_share0(d3_P2_25_s0), .output_share1(d3_P2_25_s1));
  reg_module u_reg_P2_26_d3 (.clk(clk), .input_share0(d2_P2_26_s0), .input_share1(d2_P2_26_s1), .output_share0(d3_P2_26_s0), .output_share1(d3_P2_26_s1));
  reg_module u_reg_P2_27_d3 (.clk(clk), .input_share0(d2_P2_27_s0), .input_share1(d2_P2_27_s1), .output_share0(d3_P2_27_s0), .output_share1(d3_P2_27_s1));
  reg_module u_reg_P2_28_d3 (.clk(clk), .input_share0(d2_P2_28_s0), .input_share1(d2_P2_28_s1), .output_share0(d3_P2_28_s0), .output_share1(d3_P2_28_s1));
  reg_module u_reg_P2_29_d3 (.clk(clk), .input_share0(d2_P2_29_s0), .input_share1(d2_P2_29_s1), .output_share0(d3_P2_29_s0), .output_share1(d3_P2_29_s1));
  reg_module u_reg_P2_30_d3 (.clk(clk), .input_share0(d2_P2_30_s0), .input_share1(d2_P2_30_s1), .output_share0(d3_P2_30_s0), .output_share1(d3_P2_30_s1));
  reg_module u_reg_P2_31_d3 (.clk(clk), .input_share0(d2_P2_31_s0), .input_share1(d2_P2_31_s1), .output_share0(d3_P2_31_s0), .output_share1(d3_P2_31_s1));
  reg_module u_reg_P2_7_d3 (.clk(clk), .input_share0(d2_P2_7_s0), .input_share1(d2_P2_7_s1), .output_share0(d3_P2_7_s0), .output_share1(d3_P2_7_s1));
  reg_module u_reg_P2_8_d3 (.clk(clk), .input_share0(d2_P2_8_s0), .input_share1(d2_P2_8_s1), .output_share0(d3_P2_8_s0), .output_share1(d3_P2_8_s1));
  reg_module u_reg_P2_9_d3 (.clk(clk), .input_share0(d2_P2_9_s0), .input_share1(d2_P2_9_s1), .output_share0(d3_P2_9_s0), .output_share1(d3_P2_9_s1));
  xor_module u_xor_G2_10_d3 (.x_share0(d3_t39_s0), .x_share1(d3_t39_s1), .y_share0(d3_G1_10_s0), .y_share1(d3_G1_10_s1), .z_share0(d3_G2_10_s0), .z_share1(d3_G2_10_s1));
  xor_module u_xor_G2_11_d3 (.x_share0(d3_t40_s0), .x_share1(d3_t40_s1), .y_share0(d3_G1_11_s0), .y_share1(d3_G1_11_s1), .z_share0(d3_G2_11_s0), .z_share1(d3_G2_11_s1));
  xor_module u_xor_G2_12_d3 (.x_share0(d3_t41_s0), .x_share1(d3_t41_s1), .y_share0(d3_G1_12_s0), .y_share1(d3_G1_12_s1), .z_share0(d3_G2_12_s0), .z_share1(d3_G2_12_s1));
  xor_module u_xor_G2_13_d3 (.x_share0(d3_t42_s0), .x_share1(d3_t42_s1), .y_share0(d3_G1_13_s0), .y_share1(d3_G1_13_s1), .z_share0(d3_G2_13_s0), .z_share1(d3_G2_13_s1));
  xor_module u_xor_G2_14_d3 (.x_share0(d3_t43_s0), .x_share1(d3_t43_s1), .y_share0(d3_G1_14_s0), .y_share1(d3_G1_14_s1), .z_share0(d3_G2_14_s0), .z_share1(d3_G2_14_s1));
  xor_module u_xor_G2_15_d3 (.x_share0(d3_t44_s0), .x_share1(d3_t44_s1), .y_share0(d3_G1_15_s0), .y_share1(d3_G1_15_s1), .z_share0(d3_G2_15_s0), .z_share1(d3_G2_15_s1));
  xor_module u_xor_G2_16_d3 (.x_share0(d3_t45_s0), .x_share1(d3_t45_s1), .y_share0(d3_G1_16_s0), .y_share1(d3_G1_16_s1), .z_share0(d3_G2_16_s0), .z_share1(d3_G2_16_s1));
  xor_module u_xor_G2_17_d3 (.x_share0(d3_t46_s0), .x_share1(d3_t46_s1), .y_share0(d3_G1_17_s0), .y_share1(d3_G1_17_s1), .z_share0(d3_G2_17_s0), .z_share1(d3_G2_17_s1));
  xor_module u_xor_G2_18_d3 (.x_share0(d3_t47_s0), .x_share1(d3_t47_s1), .y_share0(d3_G1_18_s0), .y_share1(d3_G1_18_s1), .z_share0(d3_G2_18_s0), .z_share1(d3_G2_18_s1));
  xor_module u_xor_G2_19_d3 (.x_share0(d3_t48_s0), .x_share1(d3_t48_s1), .y_share0(d3_G1_19_s0), .y_share1(d3_G1_19_s1), .z_share0(d3_G2_19_s0), .z_share1(d3_G2_19_s1));
  xor_module u_xor_G2_20_d3 (.x_share0(d3_t49_s0), .x_share1(d3_t49_s1), .y_share0(d3_G1_20_s0), .y_share1(d3_G1_20_s1), .z_share0(d3_G2_20_s0), .z_share1(d3_G2_20_s1));
  xor_module u_xor_G2_21_d3 (.x_share0(d3_t50_s0), .x_share1(d3_t50_s1), .y_share0(d3_G1_21_s0), .y_share1(d3_G1_21_s1), .z_share0(d3_G2_21_s0), .z_share1(d3_G2_21_s1));
  xor_module u_xor_G2_22_d3 (.x_share0(d3_t51_s0), .x_share1(d3_t51_s1), .y_share0(d3_G1_22_s0), .y_share1(d3_G1_22_s1), .z_share0(d3_G2_22_s0), .z_share1(d3_G2_22_s1));
  xor_module u_xor_G2_23_d3 (.x_share0(d3_t52_s0), .x_share1(d3_t52_s1), .y_share0(d3_G1_23_s0), .y_share1(d3_G1_23_s1), .z_share0(d3_G2_23_s0), .z_share1(d3_G2_23_s1));
  xor_module u_xor_G2_24_d3 (.x_share0(d3_t53_s0), .x_share1(d3_t53_s1), .y_share0(d3_G1_24_s0), .y_share1(d3_G1_24_s1), .z_share0(d3_G2_24_s0), .z_share1(d3_G2_24_s1));
  xor_module u_xor_G2_25_d3 (.x_share0(d3_t54_s0), .x_share1(d3_t54_s1), .y_share0(d3_G1_25_s0), .y_share1(d3_G1_25_s1), .z_share0(d3_G2_25_s0), .z_share1(d3_G2_25_s1));
  xor_module u_xor_G2_26_d3 (.x_share0(d3_t55_s0), .x_share1(d3_t55_s1), .y_share0(d3_G1_26_s0), .y_share1(d3_G1_26_s1), .z_share0(d3_G2_26_s0), .z_share1(d3_G2_26_s1));
  xor_module u_xor_G2_27_d3 (.x_share0(d3_t56_s0), .x_share1(d3_t56_s1), .y_share0(d3_G1_27_s0), .y_share1(d3_G1_27_s1), .z_share0(d3_G2_27_s0), .z_share1(d3_G2_27_s1));
  xor_module u_xor_G2_28_d3 (.x_share0(d3_t57_s0), .x_share1(d3_t57_s1), .y_share0(d3_G1_28_s0), .y_share1(d3_G1_28_s1), .z_share0(d3_G2_28_s0), .z_share1(d3_G2_28_s1));
  xor_module u_xor_G2_29_d3 (.x_share0(d3_t58_s0), .x_share1(d3_t58_s1), .y_share0(d3_G1_29_s0), .y_share1(d3_G1_29_s1), .z_share0(d3_G2_29_s0), .z_share1(d3_G2_29_s1));
  xor_module u_xor_G2_3_d3 (.x_share0(d3_t32_s0), .x_share1(d3_t32_s1), .y_share0(d3_G1_3_s0), .y_share1(d3_G1_3_s1), .z_share0(d3_G2_3_s0), .z_share1(d3_G2_3_s1));
  xor_module u_xor_G2_30_d3 (.x_share0(d3_t59_s0), .x_share1(d3_t59_s1), .y_share0(d3_G1_30_s0), .y_share1(d3_G1_30_s1), .z_share0(d3_G2_30_s0), .z_share1(d3_G2_30_s1));
  xor_module u_xor_G2_31_d3 (.x_share0(d3_t60_s0), .x_share1(d3_t60_s1), .y_share0(d3_G1_31_s0), .y_share1(d3_G1_31_s1), .z_share0(d3_G2_31_s0), .z_share1(d3_G2_31_s1));
  xor_module u_xor_G2_4_d3 (.x_share0(d3_t33_s0), .x_share1(d3_t33_s1), .y_share0(d3_G1_4_s0), .y_share1(d3_G1_4_s1), .z_share0(d3_G2_4_s0), .z_share1(d3_G2_4_s1));
  xor_module u_xor_G2_5_d3 (.x_share0(d3_t34_s0), .x_share1(d3_t34_s1), .y_share0(d3_G1_5_s0), .y_share1(d3_G1_5_s1), .z_share0(d3_G2_5_s0), .z_share1(d3_G2_5_s1));
  xor_module u_xor_G2_6_d3 (.x_share0(d3_t35_s0), .x_share1(d3_t35_s1), .y_share0(d3_G1_6_s0), .y_share1(d3_G1_6_s1), .z_share0(d3_G2_6_s0), .z_share1(d3_G2_6_s1));
  xor_module u_xor_G2_7_d3 (.x_share0(d3_t36_s0), .x_share1(d3_t36_s1), .y_share0(d3_G1_7_s0), .y_share1(d3_G1_7_s1), .z_share0(d3_G2_7_s0), .z_share1(d3_G2_7_s1));
  xor_module u_xor_G2_8_d3 (.x_share0(d3_t37_s0), .x_share1(d3_t37_s1), .y_share0(d3_G1_8_s0), .y_share1(d3_G1_8_s1), .z_share0(d3_G2_8_s0), .z_share1(d3_G2_8_s1));
  xor_module u_xor_G2_9_d3 (.x_share0(d3_t38_s0), .x_share1(d3_t38_s1), .y_share0(d3_G1_9_s0), .y_share1(d3_G1_9_s1), .z_share0(d3_G2_9_s0), .z_share1(d3_G2_9_s1));
  xor_module u_xor_G3_4_d3 (.x_share0(d3_t61_s0), .x_share1(d3_t61_s1), .y_share0(d3_G2_4_s0), .y_share1(d3_G2_4_s1), .z_share0(d3_G3_4_s0), .z_share1(d3_G3_4_s1));
  xor_module u_xor_G3_5_d3 (.x_share0(d3_t62_s0), .x_share1(d3_t62_s1), .y_share0(d3_G2_5_s0), .y_share1(d3_G2_5_s1), .z_share0(d3_G3_5_s0), .z_share1(d3_G3_5_s1));
  xor_module u_xor_G3_6_d3 (.x_share0(d3_t63_s0), .x_share1(d3_t63_s1), .y_share0(d3_G2_6_s0), .y_share1(d3_G2_6_s1), .z_share0(d3_G3_6_s0), .z_share1(d3_G3_6_s1));
  and_module u_and_P3_10_d3 (.clk(clk), .x_share0(d2_P2_10_s0), .x_share1(d2_P2_10_s1), .y_share0(d2_P2_6_s0), .y_share1(d2_P2_6_s1), .rand(r_P3_10), .z_share0(d3_P3_10_s0), .z_share1(d3_P3_10_s1));
  assign r_P3_10 = stage3_share0[22];
  and_module u_and_P3_11_d3 (.clk(clk), .x_share0(d2_P2_11_s0), .x_share1(d2_P2_11_s1), .y_share0(d2_P2_7_s0), .y_share1(d2_P2_7_s1), .rand(r_P3_11), .z_share0(d3_P3_11_s0), .z_share1(d3_P3_11_s1));
  assign r_P3_11 = stage3_share0[6];
  and_module u_and_P3_12_d3 (.clk(clk), .x_share0(d2_P2_12_s0), .x_share1(d2_P2_12_s1), .y_share0(d2_P2_8_s0), .y_share1(d2_P2_8_s1), .rand(r_P3_12), .z_share0(d3_P3_12_s0), .z_share1(d3_P3_12_s1));
  assign r_P3_12 = stage3_share0[18];
  and_module u_and_P3_13_d3 (.clk(clk), .x_share0(d2_P2_13_s0), .x_share1(d2_P2_13_s1), .y_share0(d2_P2_9_s0), .y_share1(d2_P2_9_s1), .rand(r_P3_13), .z_share0(d3_P3_13_s0), .z_share1(d3_P3_13_s1));
  assign r_P3_13 = stage3_share0[18];
  and_module u_and_P3_14_d3 (.clk(clk), .x_share0(d2_P2_14_s0), .x_share1(d2_P2_14_s1), .y_share0(d2_P2_10_s0), .y_share1(d2_P2_10_s1), .rand(r_P3_14), .z_share0(d3_P3_14_s0), .z_share1(d3_P3_14_s1));
  assign r_P3_14 = stage3_share0[9];
  and_module u_and_P3_15_d3 (.clk(clk), .x_share0(d2_P2_15_s0), .x_share1(d2_P2_15_s1), .y_share0(d2_P2_11_s0), .y_share1(d2_P2_11_s1), .rand(r_P3_15), .z_share0(d3_P3_15_s0), .z_share1(d3_P3_15_s1));
  assign r_P3_15 = stage3_share0[3];
  and_module u_and_P3_16_d3 (.clk(clk), .x_share0(d2_P2_16_s0), .x_share1(d2_P2_16_s1), .y_share0(d2_P2_12_s0), .y_share1(d2_P2_12_s1), .rand(r_P3_16), .z_share0(d3_P3_16_s0), .z_share1(d3_P3_16_s1));
  assign r_P3_16 = stage3_share0[10];
  and_module u_and_P3_17_d3 (.clk(clk), .x_share0(d2_P2_17_s0), .x_share1(d2_P2_17_s1), .y_share0(d2_P2_13_s0), .y_share1(d2_P2_13_s1), .rand(r_P3_17), .z_share0(d3_P3_17_s0), .z_share1(d3_P3_17_s1));
  assign r_P3_17 = stage3_share0[20];
  and_module u_and_P3_18_d3 (.clk(clk), .x_share0(d2_P2_18_s0), .x_share1(d2_P2_18_s1), .y_share0(d2_P2_14_s0), .y_share1(d2_P2_14_s1), .rand(r_P3_18), .z_share0(d3_P3_18_s0), .z_share1(d3_P3_18_s1));
  assign r_P3_18 = stage3_share0[9];
  and_module u_and_P3_19_d3 (.clk(clk), .x_share0(d2_P2_19_s0), .x_share1(d2_P2_19_s1), .y_share0(d2_P2_15_s0), .y_share1(d2_P2_15_s1), .rand(r_P3_19), .z_share0(d3_P3_19_s0), .z_share1(d3_P3_19_s1));
  assign r_P3_19 = stage3_share0[22];
  and_module u_and_P3_20_d3 (.clk(clk), .x_share0(d2_P2_20_s0), .x_share1(d2_P2_20_s1), .y_share0(d2_P2_16_s0), .y_share1(d2_P2_16_s1), .rand(r_P3_20), .z_share0(d3_P3_20_s0), .z_share1(d3_P3_20_s1));
  assign r_P3_20 = stage3_share0[21];
  and_module u_and_P3_21_d3 (.clk(clk), .x_share0(d2_P2_21_s0), .x_share1(d2_P2_21_s1), .y_share0(d2_P2_17_s0), .y_share1(d2_P2_17_s1), .rand(r_P3_21), .z_share0(d3_P3_21_s0), .z_share1(d3_P3_21_s1));
  assign r_P3_21 = stage3_share0[23];
  and_module u_and_P3_22_d3 (.clk(clk), .x_share0(d2_P2_22_s0), .x_share1(d2_P2_22_s1), .y_share0(d2_P2_18_s0), .y_share1(d2_P2_18_s1), .rand(r_P3_22), .z_share0(d3_P3_22_s0), .z_share1(d3_P3_22_s1));
  assign r_P3_22 = stage3_share0[23];
  and_module u_and_P3_23_d3 (.clk(clk), .x_share0(d2_P2_23_s0), .x_share1(d2_P2_23_s1), .y_share0(d2_P2_19_s0), .y_share1(d2_P2_19_s1), .rand(r_P3_23), .z_share0(d3_P3_23_s0), .z_share1(d3_P3_23_s1));
  assign r_P3_23 = stage3_share0[17];
  and_module u_and_P3_24_d3 (.clk(clk), .x_share0(d2_P2_24_s0), .x_share1(d2_P2_24_s1), .y_share0(d2_P2_20_s0), .y_share1(d2_P2_20_s1), .rand(r_P3_24), .z_share0(d3_P3_24_s0), .z_share1(d3_P3_24_s1));
  assign r_P3_24 = stage3_share0[8];
  and_module u_and_P3_25_d3 (.clk(clk), .x_share0(d2_P2_25_s0), .x_share1(d2_P2_25_s1), .y_share0(d2_P2_21_s0), .y_share1(d2_P2_21_s1), .rand(r_P3_25), .z_share0(d3_P3_25_s0), .z_share1(d3_P3_25_s1));
  assign r_P3_25 = stage3_share0[4];
  and_module u_and_P3_26_d3 (.clk(clk), .x_share0(d2_P2_26_s0), .x_share1(d2_P2_26_s1), .y_share0(d2_P2_22_s0), .y_share1(d2_P2_22_s1), .rand(r_P3_26), .z_share0(d3_P3_26_s0), .z_share1(d3_P3_26_s1));
  assign r_P3_26 = stage3_share0[18];
  and_module u_and_P3_27_d3 (.clk(clk), .x_share0(d2_P2_27_s0), .x_share1(d2_P2_27_s1), .y_share0(d2_P2_23_s0), .y_share1(d2_P2_23_s1), .rand(r_P3_27), .z_share0(d3_P3_27_s0), .z_share1(d3_P3_27_s1));
  assign r_P3_27 = stage3_share0[17];
  and_module u_and_P3_28_d3 (.clk(clk), .x_share0(d2_P2_28_s0), .x_share1(d2_P2_28_s1), .y_share0(d2_P2_24_s0), .y_share1(d2_P2_24_s1), .rand(r_P3_28), .z_share0(d3_P3_28_s0), .z_share1(d3_P3_28_s1));
  assign r_P3_28 = stage3_share0[20];
  and_module u_and_P3_29_d3 (.clk(clk), .x_share0(d2_P2_29_s0), .x_share1(d2_P2_29_s1), .y_share0(d2_P2_25_s0), .y_share1(d2_P2_25_s1), .rand(r_P3_29), .z_share0(d3_P3_29_s0), .z_share1(d3_P3_29_s1));
  assign r_P3_29 = stage3_share0[22];
  and_module u_and_P3_30_d3 (.clk(clk), .x_share0(d2_P2_30_s0), .x_share1(d2_P2_30_s1), .y_share0(d2_P2_26_s0), .y_share1(d2_P2_26_s1), .rand(r_P3_30), .z_share0(d3_P3_30_s0), .z_share1(d3_P3_30_s1));
  assign r_P3_30 = stage3_share0[22];
  and_module u_and_P3_31_d3 (.clk(clk), .x_share0(d2_P2_31_s0), .x_share1(d2_P2_31_s1), .y_share0(d2_P2_27_s0), .y_share1(d2_P2_27_s1), .rand(r_P3_31), .z_share0(d3_P3_31_s0), .z_share1(d3_P3_31_s1));
  assign r_P3_31 = stage3_share0[21];
  and_module u_and_P3_8_d3 (.clk(clk), .x_share0(d2_P2_8_s0), .x_share1(d2_P2_8_s1), .y_share0(d2_P2_4_s0), .y_share1(d2_P2_4_s1), .rand(r_P3_8), .z_share0(d3_P3_8_s0), .z_share1(d3_P3_8_s1));
  assign r_P3_8 = stage3_share0[17];
  and_module u_and_P3_9_d3 (.clk(clk), .x_share0(d2_P2_9_s0), .x_share1(d2_P2_9_s1), .y_share0(d2_P2_5_s0), .y_share1(d2_P2_5_s1), .rand(r_P3_9), .z_share0(d3_P3_9_s0), .z_share1(d3_P3_9_s1));
  assign r_P3_9 = stage3_share0[7];
  xor_module u_xor_o4_d3 (.x_share0(d3_P0_4_s0), .x_share1(d3_P0_4_s1), .y_share0(d3_G2_3_s0), .y_share1(d3_G2_3_s1), .z_share0(d3_o4_s0), .z_share1(d3_o4_s1));
  xor_module u_xor_o5_d3 (.x_share0(d3_P0_5_s0), .x_share1(d3_P0_5_s1), .y_share0(d3_G3_4_s0), .y_share1(d3_G3_4_s1), .z_share0(d3_o5_s0), .z_share1(d3_o5_s1));
  xor_module u_xor_o6_d3 (.x_share0(d3_P0_6_s0), .x_share1(d3_P0_6_s1), .y_share0(d3_G3_5_s0), .y_share1(d3_G3_5_s1), .z_share0(d3_o6_s0), .z_share1(d3_o6_s1));
  xor_module u_xor_o7_d3 (.x_share0(d3_P0_7_s0), .x_share1(d3_P0_7_s1), .y_share0(d3_G3_6_s0), .y_share1(d3_G3_6_s1), .z_share0(d3_o7_s0), .z_share1(d3_o7_s1));
  and_module u_and_t32_d3 (.clk(clk), .x_share0(d2_P1_3_s0), .x_share1(d2_P1_3_s1), .y_share0(d2_G1_1_s0), .y_share1(d2_G1_1_s1), .rand(r_t32), .z_share0(d3_t32_s0), .z_share1(d3_t32_s1));
  assign r_t32 = stage3_share0[21];
  and_module u_and_t33_d3 (.clk(clk), .x_share0(d2_P1_4_s0), .x_share1(d2_P1_4_s1), .y_share0(d2_G1_2_s0), .y_share1(d2_G1_2_s1), .rand(r_t33), .z_share0(d3_t33_s0), .z_share1(d3_t33_s1));
  assign r_t33 = stage3_share0[15];
  and_module u_and_t34_d3 (.clk(clk), .x_share0(d2_P1_5_s0), .x_share1(d2_P1_5_s1), .y_share0(d2_G1_3_s0), .y_share1(d2_G1_3_s1), .rand(r_t34), .z_share0(d3_t34_s0), .z_share1(d3_t34_s1));
  assign r_t34 = stage3_share0[19];
  and_module u_and_t35_d3 (.clk(clk), .x_share0(d2_P1_6_s0), .x_share1(d2_P1_6_s1), .y_share0(d2_G1_4_s0), .y_share1(d2_G1_4_s1), .rand(r_t35), .z_share0(d3_t35_s0), .z_share1(d3_t35_s1));
  assign r_t35 = stage3_share0[16];
  and_module u_and_t36_d3 (.clk(clk), .x_share0(d2_P1_7_s0), .x_share1(d2_P1_7_s1), .y_share0(d2_G1_5_s0), .y_share1(d2_G1_5_s1), .rand(r_t36), .z_share0(d3_t36_s0), .z_share1(d3_t36_s1));
  assign r_t36 = stage3_share0[19];
  and_module u_and_t37_d3 (.clk(clk), .x_share0(d2_P1_8_s0), .x_share1(d2_P1_8_s1), .y_share0(d2_G1_6_s0), .y_share1(d2_G1_6_s1), .rand(r_t37), .z_share0(d3_t37_s0), .z_share1(d3_t37_s1));
  assign r_t37 = stage3_share0[16];
  and_module u_and_t38_d3 (.clk(clk), .x_share0(d2_P1_9_s0), .x_share1(d2_P1_9_s1), .y_share0(d2_G1_7_s0), .y_share1(d2_G1_7_s1), .rand(r_t38), .z_share0(d3_t38_s0), .z_share1(d3_t38_s1));
  assign r_t38 = stage3_share0[12];
  and_module u_and_t39_d3 (.clk(clk), .x_share0(d2_P1_10_s0), .x_share1(d2_P1_10_s1), .y_share0(d2_G1_8_s0), .y_share1(d2_G1_8_s1), .rand(r_t39), .z_share0(d3_t39_s0), .z_share1(d3_t39_s1));
  assign r_t39 = stage3_share0[14];
  and_module u_and_t40_d3 (.clk(clk), .x_share0(d2_P1_11_s0), .x_share1(d2_P1_11_s1), .y_share0(d2_G1_9_s0), .y_share1(d2_G1_9_s1), .rand(r_t40), .z_share0(d3_t40_s0), .z_share1(d3_t40_s1));
  assign r_t40 = stage3_share0[3];
  and_module u_and_t41_d3 (.clk(clk), .x_share0(d2_P1_12_s0), .x_share1(d2_P1_12_s1), .y_share0(d2_G1_10_s0), .y_share1(d2_G1_10_s1), .rand(r_t41), .z_share0(d3_t41_s0), .z_share1(d3_t41_s1));
  assign r_t41 = stage3_share0[17];
  and_module u_and_t42_d3 (.clk(clk), .x_share0(d2_P1_13_s0), .x_share1(d2_P1_13_s1), .y_share0(d2_G1_11_s0), .y_share1(d2_G1_11_s1), .rand(r_t42), .z_share0(d3_t42_s0), .z_share1(d3_t42_s1));
  assign r_t42 = stage3_share0[20];
  and_module u_and_t43_d3 (.clk(clk), .x_share0(d2_P1_14_s0), .x_share1(d2_P1_14_s1), .y_share0(d2_G1_12_s0), .y_share1(d2_G1_12_s1), .rand(r_t43), .z_share0(d3_t43_s0), .z_share1(d3_t43_s1));
  assign r_t43 = stage3_share0[21];
  and_module u_and_t44_d3 (.clk(clk), .x_share0(d2_P1_15_s0), .x_share1(d2_P1_15_s1), .y_share0(d2_G1_13_s0), .y_share1(d2_G1_13_s1), .rand(r_t44), .z_share0(d3_t44_s0), .z_share1(d3_t44_s1));
  assign r_t44 = stage3_share0[15];
  and_module u_and_t45_d3 (.clk(clk), .x_share0(d2_P1_16_s0), .x_share1(d2_P1_16_s1), .y_share0(d2_G1_14_s0), .y_share1(d2_G1_14_s1), .rand(r_t45), .z_share0(d3_t45_s0), .z_share1(d3_t45_s1));
  assign r_t45 = stage3_share0[15];
  and_module u_and_t46_d3 (.clk(clk), .x_share0(d2_P1_17_s0), .x_share1(d2_P1_17_s1), .y_share0(d2_G1_15_s0), .y_share1(d2_G1_15_s1), .rand(r_t46), .z_share0(d3_t46_s0), .z_share1(d3_t46_s1));
  assign r_t46 = stage3_share0[13];
  and_module u_and_t47_d3 (.clk(clk), .x_share0(d2_P1_18_s0), .x_share1(d2_P1_18_s1), .y_share0(d2_G1_16_s0), .y_share1(d2_G1_16_s1), .rand(r_t47), .z_share0(d3_t47_s0), .z_share1(d3_t47_s1));
  assign r_t47 = stage3_share0[13];
  and_module u_and_t48_d3 (.clk(clk), .x_share0(d2_P1_19_s0), .x_share1(d2_P1_19_s1), .y_share0(d2_G1_17_s0), .y_share1(d2_G1_17_s1), .rand(r_t48), .z_share0(d3_t48_s0), .z_share1(d3_t48_s1));
  assign r_t48 = stage3_share0[16];
  and_module u_and_t49_d3 (.clk(clk), .x_share0(d2_P1_20_s0), .x_share1(d2_P1_20_s1), .y_share0(d2_G1_18_s0), .y_share1(d2_G1_18_s1), .rand(r_t49), .z_share0(d3_t49_s0), .z_share1(d3_t49_s1));
  assign r_t49 = stage3_share0[12];
  and_module u_and_t50_d3 (.clk(clk), .x_share0(d2_P1_21_s0), .x_share1(d2_P1_21_s1), .y_share0(d2_G1_19_s0), .y_share1(d2_G1_19_s1), .rand(r_t50), .z_share0(d3_t50_s0), .z_share1(d3_t50_s1));
  assign r_t50 = stage3_share0[9];
  and_module u_and_t51_d3 (.clk(clk), .x_share0(d2_P1_22_s0), .x_share1(d2_P1_22_s1), .y_share0(d2_G1_20_s0), .y_share1(d2_G1_20_s1), .rand(r_t51), .z_share0(d3_t51_s0), .z_share1(d3_t51_s1));
  assign r_t51 = stage3_share0[6];
  and_module u_and_t52_d3 (.clk(clk), .x_share0(d2_P1_23_s0), .x_share1(d2_P1_23_s1), .y_share0(d2_G1_21_s0), .y_share1(d2_G1_21_s1), .rand(r_t52), .z_share0(d3_t52_s0), .z_share1(d3_t52_s1));
  assign r_t52 = stage3_share0[13];
  and_module u_and_t53_d3 (.clk(clk), .x_share0(d2_P1_24_s0), .x_share1(d2_P1_24_s1), .y_share0(d2_G1_22_s0), .y_share1(d2_G1_22_s1), .rand(r_t53), .z_share0(d3_t53_s0), .z_share1(d3_t53_s1));
  assign r_t53 = stage3_share0[10];
  and_module u_and_t54_d3 (.clk(clk), .x_share0(d2_P1_25_s0), .x_share1(d2_P1_25_s1), .y_share0(d2_G1_23_s0), .y_share1(d2_G1_23_s1), .rand(r_t54), .z_share0(d3_t54_s0), .z_share1(d3_t54_s1));
  assign r_t54 = stage3_share0[20];
  and_module u_and_t55_d3 (.clk(clk), .x_share0(d2_P1_26_s0), .x_share1(d2_P1_26_s1), .y_share0(d2_G1_24_s0), .y_share1(d2_G1_24_s1), .rand(r_t55), .z_share0(d3_t55_s0), .z_share1(d3_t55_s1));
  assign r_t55 = stage3_share0[20];
  and_module u_and_t56_d3 (.clk(clk), .x_share0(d2_P1_27_s0), .x_share1(d2_P1_27_s1), .y_share0(d2_G1_25_s0), .y_share1(d2_G1_25_s1), .rand(r_t56), .z_share0(d3_t56_s0), .z_share1(d3_t56_s1));
  assign r_t56 = stage3_share0[4];
  and_module u_and_t57_d3 (.clk(clk), .x_share0(d2_P1_28_s0), .x_share1(d2_P1_28_s1), .y_share0(d2_G1_26_s0), .y_share1(d2_G1_26_s1), .rand(r_t57), .z_share0(d3_t57_s0), .z_share1(d3_t57_s1));
  assign r_t57 = stage3_share0[15];
  and_module u_and_t58_d3 (.clk(clk), .x_share0(d2_P1_29_s0), .x_share1(d2_P1_29_s1), .y_share0(d2_G1_27_s0), .y_share1(d2_G1_27_s1), .rand(r_t58), .z_share0(d3_t58_s0), .z_share1(d3_t58_s1));
  assign r_t58 = stage3_share0[13];
  and_module u_and_t59_d3 (.clk(clk), .x_share0(d2_P1_30_s0), .x_share1(d2_P1_30_s1), .y_share0(d2_G1_28_s0), .y_share1(d2_G1_28_s1), .rand(r_t59), .z_share0(d3_t59_s0), .z_share1(d3_t59_s1));
  assign r_t59 = stage3_share0[11];
  and_module u_and_t60_d3 (.clk(clk), .x_share0(d2_P1_31_s0), .x_share1(d2_P1_31_s1), .y_share0(d2_G1_29_s0), .y_share1(d2_G1_29_s1), .rand(r_t60), .z_share0(d3_t60_s0), .z_share1(d3_t60_s1));
  assign r_t60 = stage3_share0[17];
  and_module u_and_t61_d3 (.clk(clk), .x_share0(d2_P2_4_s0), .x_share1(d2_P2_4_s1), .y_share0(d2_G0_0_s0), .y_share1(d2_G0_0_s1), .rand(r_t61), .z_share0(d3_t61_s0), .z_share1(d3_t61_s1));
  assign r_t61 = stage3_share0[24];
  and_module u_and_t62_d3 (.clk(clk), .x_share0(d2_P2_5_s0), .x_share1(d2_P2_5_s1), .y_share0(d2_G1_1_s0), .y_share1(d2_G1_1_s1), .rand(r_t62), .z_share0(d3_t62_s0), .z_share1(d3_t62_s1));
  assign r_t62 = stage3_share0[16];
  and_module u_and_t63_d3 (.clk(clk), .x_share0(d2_P2_6_s0), .x_share1(d2_P2_6_s1), .y_share0(d2_G2_2_s0), .y_share1(d2_G2_2_s1), .rand(r_t63), .z_share0(d3_t63_s0), .z_share1(d3_t63_s1));
  assign r_t63 = stage3_share0[3];
  reg_module u_reg_G0_0_d4 (.clk(clk), .input_share0(d3_G0_0_s0), .input_share1(d3_G0_0_s1), .output_share0(d4_G0_0_s0), .output_share1(d4_G0_0_s1));
  reg_module u_reg_G1_1_d4 (.clk(clk), .input_share0(d3_G1_1_s0), .input_share1(d3_G1_1_s1), .output_share0(d4_G1_1_s0), .output_share1(d4_G1_1_s1));
  reg_module u_reg_G2_10_d4 (.clk(clk), .input_share0(d3_G2_10_s0), .input_share1(d3_G2_10_s1), .output_share0(d4_G2_10_s0), .output_share1(d4_G2_10_s1));
  reg_module u_reg_G2_11_d4 (.clk(clk), .input_share0(d3_G2_11_s0), .input_share1(d3_G2_11_s1), .output_share0(d4_G2_11_s0), .output_share1(d4_G2_11_s1));
  reg_module u_reg_G2_12_d4 (.clk(clk), .input_share0(d3_G2_12_s0), .input_share1(d3_G2_12_s1), .output_share0(d4_G2_12_s0), .output_share1(d4_G2_12_s1));
  reg_module u_reg_G2_13_d4 (.clk(clk), .input_share0(d3_G2_13_s0), .input_share1(d3_G2_13_s1), .output_share0(d4_G2_13_s0), .output_share1(d4_G2_13_s1));
  reg_module u_reg_G2_14_d4 (.clk(clk), .input_share0(d3_G2_14_s0), .input_share1(d3_G2_14_s1), .output_share0(d4_G2_14_s0), .output_share1(d4_G2_14_s1));
  reg_module u_reg_G2_15_d4 (.clk(clk), .input_share0(d3_G2_15_s0), .input_share1(d3_G2_15_s1), .output_share0(d4_G2_15_s0), .output_share1(d4_G2_15_s1));
  reg_module u_reg_G2_16_d4 (.clk(clk), .input_share0(d3_G2_16_s0), .input_share1(d3_G2_16_s1), .output_share0(d4_G2_16_s0), .output_share1(d4_G2_16_s1));
  reg_module u_reg_G2_17_d4 (.clk(clk), .input_share0(d3_G2_17_s0), .input_share1(d3_G2_17_s1), .output_share0(d4_G2_17_s0), .output_share1(d4_G2_17_s1));
  reg_module u_reg_G2_18_d4 (.clk(clk), .input_share0(d3_G2_18_s0), .input_share1(d3_G2_18_s1), .output_share0(d4_G2_18_s0), .output_share1(d4_G2_18_s1));
  reg_module u_reg_G2_19_d4 (.clk(clk), .input_share0(d3_G2_19_s0), .input_share1(d3_G2_19_s1), .output_share0(d4_G2_19_s0), .output_share1(d4_G2_19_s1));
  reg_module u_reg_G2_2_d4 (.clk(clk), .input_share0(d3_G2_2_s0), .input_share1(d3_G2_2_s1), .output_share0(d4_G2_2_s0), .output_share1(d4_G2_2_s1));
  reg_module u_reg_G2_20_d4 (.clk(clk), .input_share0(d3_G2_20_s0), .input_share1(d3_G2_20_s1), .output_share0(d4_G2_20_s0), .output_share1(d4_G2_20_s1));
  reg_module u_reg_G2_21_d4 (.clk(clk), .input_share0(d3_G2_21_s0), .input_share1(d3_G2_21_s1), .output_share0(d4_G2_21_s0), .output_share1(d4_G2_21_s1));
  reg_module u_reg_G2_22_d4 (.clk(clk), .input_share0(d3_G2_22_s0), .input_share1(d3_G2_22_s1), .output_share0(d4_G2_22_s0), .output_share1(d4_G2_22_s1));
  reg_module u_reg_G2_23_d4 (.clk(clk), .input_share0(d3_G2_23_s0), .input_share1(d3_G2_23_s1), .output_share0(d4_G2_23_s0), .output_share1(d4_G2_23_s1));
  reg_module u_reg_G2_24_d4 (.clk(clk), .input_share0(d3_G2_24_s0), .input_share1(d3_G2_24_s1), .output_share0(d4_G2_24_s0), .output_share1(d4_G2_24_s1));
  reg_module u_reg_G2_25_d4 (.clk(clk), .input_share0(d3_G2_25_s0), .input_share1(d3_G2_25_s1), .output_share0(d4_G2_25_s0), .output_share1(d4_G2_25_s1));
  reg_module u_reg_G2_26_d4 (.clk(clk), .input_share0(d3_G2_26_s0), .input_share1(d3_G2_26_s1), .output_share0(d4_G2_26_s0), .output_share1(d4_G2_26_s1));
  reg_module u_reg_G2_27_d4 (.clk(clk), .input_share0(d3_G2_27_s0), .input_share1(d3_G2_27_s1), .output_share0(d4_G2_27_s0), .output_share1(d4_G2_27_s1));
  reg_module u_reg_G2_28_d4 (.clk(clk), .input_share0(d3_G2_28_s0), .input_share1(d3_G2_28_s1), .output_share0(d4_G2_28_s0), .output_share1(d4_G2_28_s1));
  reg_module u_reg_G2_29_d4 (.clk(clk), .input_share0(d3_G2_29_s0), .input_share1(d3_G2_29_s1), .output_share0(d4_G2_29_s0), .output_share1(d4_G2_29_s1));
  reg_module u_reg_G2_3_d4 (.clk(clk), .input_share0(d3_G2_3_s0), .input_share1(d3_G2_3_s1), .output_share0(d4_G2_3_s0), .output_share1(d4_G2_3_s1));
  reg_module u_reg_G2_30_d4 (.clk(clk), .input_share0(d3_G2_30_s0), .input_share1(d3_G2_30_s1), .output_share0(d4_G2_30_s0), .output_share1(d4_G2_30_s1));
  reg_module u_reg_G2_31_d4 (.clk(clk), .input_share0(d3_G2_31_s0), .input_share1(d3_G2_31_s1), .output_share0(d4_G2_31_s0), .output_share1(d4_G2_31_s1));
  reg_module u_reg_G2_7_d4 (.clk(clk), .input_share0(d3_G2_7_s0), .input_share1(d3_G2_7_s1), .output_share0(d4_G2_7_s0), .output_share1(d4_G2_7_s1));
  reg_module u_reg_G2_8_d4 (.clk(clk), .input_share0(d3_G2_8_s0), .input_share1(d3_G2_8_s1), .output_share0(d4_G2_8_s0), .output_share1(d4_G2_8_s1));
  reg_module u_reg_G2_9_d4 (.clk(clk), .input_share0(d3_G2_9_s0), .input_share1(d3_G2_9_s1), .output_share0(d4_G2_9_s0), .output_share1(d4_G2_9_s1));
  reg_module u_reg_G3_4_d4 (.clk(clk), .input_share0(d3_G3_4_s0), .input_share1(d3_G3_4_s1), .output_share0(d4_G3_4_s0), .output_share1(d4_G3_4_s1));
  reg_module u_reg_G3_5_d4 (.clk(clk), .input_share0(d3_G3_5_s0), .input_share1(d3_G3_5_s1), .output_share0(d4_G3_5_s0), .output_share1(d4_G3_5_s1));
  reg_module u_reg_G3_6_d4 (.clk(clk), .input_share0(d3_G3_6_s0), .input_share1(d3_G3_6_s1), .output_share0(d4_G3_6_s0), .output_share1(d4_G3_6_s1));
  reg_module u_reg_P0_10_d4 (.clk(clk), .input_share0(d3_P0_10_s0), .input_share1(d3_P0_10_s1), .output_share0(d4_P0_10_s0), .output_share1(d4_P0_10_s1));
  reg_module u_reg_P0_11_d4 (.clk(clk), .input_share0(d3_P0_11_s0), .input_share1(d3_P0_11_s1), .output_share0(d4_P0_11_s0), .output_share1(d4_P0_11_s1));
  reg_module u_reg_P0_12_d4 (.clk(clk), .input_share0(d3_P0_12_s0), .input_share1(d3_P0_12_s1), .output_share0(d4_P0_12_s0), .output_share1(d4_P0_12_s1));
  reg_module u_reg_P0_13_d4 (.clk(clk), .input_share0(d3_P0_13_s0), .input_share1(d3_P0_13_s1), .output_share0(d4_P0_13_s0), .output_share1(d4_P0_13_s1));
  reg_module u_reg_P0_14_d4 (.clk(clk), .input_share0(d3_P0_14_s0), .input_share1(d3_P0_14_s1), .output_share0(d4_P0_14_s0), .output_share1(d4_P0_14_s1));
  reg_module u_reg_P0_15_d4 (.clk(clk), .input_share0(d3_P0_15_s0), .input_share1(d3_P0_15_s1), .output_share0(d4_P0_15_s0), .output_share1(d4_P0_15_s1));
  reg_module u_reg_P0_16_d4 (.clk(clk), .input_share0(d3_P0_16_s0), .input_share1(d3_P0_16_s1), .output_share0(d4_P0_16_s0), .output_share1(d4_P0_16_s1));
  reg_module u_reg_P0_17_d4 (.clk(clk), .input_share0(d3_P0_17_s0), .input_share1(d3_P0_17_s1), .output_share0(d4_P0_17_s0), .output_share1(d4_P0_17_s1));
  reg_module u_reg_P0_18_d4 (.clk(clk), .input_share0(d3_P0_18_s0), .input_share1(d3_P0_18_s1), .output_share0(d4_P0_18_s0), .output_share1(d4_P0_18_s1));
  reg_module u_reg_P0_19_d4 (.clk(clk), .input_share0(d3_P0_19_s0), .input_share1(d3_P0_19_s1), .output_share0(d4_P0_19_s0), .output_share1(d4_P0_19_s1));
  reg_module u_reg_P0_20_d4 (.clk(clk), .input_share0(d3_P0_20_s0), .input_share1(d3_P0_20_s1), .output_share0(d4_P0_20_s0), .output_share1(d4_P0_20_s1));
  reg_module u_reg_P0_21_d4 (.clk(clk), .input_share0(d3_P0_21_s0), .input_share1(d3_P0_21_s1), .output_share0(d4_P0_21_s0), .output_share1(d4_P0_21_s1));
  reg_module u_reg_P0_22_d4 (.clk(clk), .input_share0(d3_P0_22_s0), .input_share1(d3_P0_22_s1), .output_share0(d4_P0_22_s0), .output_share1(d4_P0_22_s1));
  reg_module u_reg_P0_23_d4 (.clk(clk), .input_share0(d3_P0_23_s0), .input_share1(d3_P0_23_s1), .output_share0(d4_P0_23_s0), .output_share1(d4_P0_23_s1));
  reg_module u_reg_P0_24_d4 (.clk(clk), .input_share0(d3_P0_24_s0), .input_share1(d3_P0_24_s1), .output_share0(d4_P0_24_s0), .output_share1(d4_P0_24_s1));
  reg_module u_reg_P0_25_d4 (.clk(clk), .input_share0(d3_P0_25_s0), .input_share1(d3_P0_25_s1), .output_share0(d4_P0_25_s0), .output_share1(d4_P0_25_s1));
  reg_module u_reg_P0_26_d4 (.clk(clk), .input_share0(d3_P0_26_s0), .input_share1(d3_P0_26_s1), .output_share0(d4_P0_26_s0), .output_share1(d4_P0_26_s1));
  reg_module u_reg_P0_27_d4 (.clk(clk), .input_share0(d3_P0_27_s0), .input_share1(d3_P0_27_s1), .output_share0(d4_P0_27_s0), .output_share1(d4_P0_27_s1));
  reg_module u_reg_P0_28_d4 (.clk(clk), .input_share0(d3_P0_28_s0), .input_share1(d3_P0_28_s1), .output_share0(d4_P0_28_s0), .output_share1(d4_P0_28_s1));
  reg_module u_reg_P0_29_d4 (.clk(clk), .input_share0(d3_P0_29_s0), .input_share1(d3_P0_29_s1), .output_share0(d4_P0_29_s0), .output_share1(d4_P0_29_s1));
  reg_module u_reg_P0_30_d4 (.clk(clk), .input_share0(d3_P0_30_s0), .input_share1(d3_P0_30_s1), .output_share0(d4_P0_30_s0), .output_share1(d4_P0_30_s1));
  reg_module u_reg_P0_31_d4 (.clk(clk), .input_share0(d3_P0_31_s0), .input_share1(d3_P0_31_s1), .output_share0(d4_P0_31_s0), .output_share1(d4_P0_31_s1));
  reg_module u_reg_P0_8_d4 (.clk(clk), .input_share0(d3_P0_8_s0), .input_share1(d3_P0_8_s1), .output_share0(d4_P0_8_s0), .output_share1(d4_P0_8_s1));
  reg_module u_reg_P0_9_d4 (.clk(clk), .input_share0(d3_P0_9_s0), .input_share1(d3_P0_9_s1), .output_share0(d4_P0_9_s0), .output_share1(d4_P0_9_s1));
  reg_module u_reg_P3_15_d4 (.clk(clk), .input_share0(d3_P3_15_s0), .input_share1(d3_P3_15_s1), .output_share0(d4_P3_15_s0), .output_share1(d4_P3_15_s1));
  reg_module u_reg_P3_16_d4 (.clk(clk), .input_share0(d3_P3_16_s0), .input_share1(d3_P3_16_s1), .output_share0(d4_P3_16_s0), .output_share1(d4_P3_16_s1));
  reg_module u_reg_P3_17_d4 (.clk(clk), .input_share0(d3_P3_17_s0), .input_share1(d3_P3_17_s1), .output_share0(d4_P3_17_s0), .output_share1(d4_P3_17_s1));
  reg_module u_reg_P3_18_d4 (.clk(clk), .input_share0(d3_P3_18_s0), .input_share1(d3_P3_18_s1), .output_share0(d4_P3_18_s0), .output_share1(d4_P3_18_s1));
  reg_module u_reg_P3_19_d4 (.clk(clk), .input_share0(d3_P3_19_s0), .input_share1(d3_P3_19_s1), .output_share0(d4_P3_19_s0), .output_share1(d4_P3_19_s1));
  reg_module u_reg_P3_20_d4 (.clk(clk), .input_share0(d3_P3_20_s0), .input_share1(d3_P3_20_s1), .output_share0(d4_P3_20_s0), .output_share1(d4_P3_20_s1));
  reg_module u_reg_P3_21_d4 (.clk(clk), .input_share0(d3_P3_21_s0), .input_share1(d3_P3_21_s1), .output_share0(d4_P3_21_s0), .output_share1(d4_P3_21_s1));
  reg_module u_reg_P3_22_d4 (.clk(clk), .input_share0(d3_P3_22_s0), .input_share1(d3_P3_22_s1), .output_share0(d4_P3_22_s0), .output_share1(d4_P3_22_s1));
  reg_module u_reg_P3_23_d4 (.clk(clk), .input_share0(d3_P3_23_s0), .input_share1(d3_P3_23_s1), .output_share0(d4_P3_23_s0), .output_share1(d4_P3_23_s1));
  reg_module u_reg_P3_24_d4 (.clk(clk), .input_share0(d3_P3_24_s0), .input_share1(d3_P3_24_s1), .output_share0(d4_P3_24_s0), .output_share1(d4_P3_24_s1));
  reg_module u_reg_P3_25_d4 (.clk(clk), .input_share0(d3_P3_25_s0), .input_share1(d3_P3_25_s1), .output_share0(d4_P3_25_s0), .output_share1(d4_P3_25_s1));
  reg_module u_reg_P3_26_d4 (.clk(clk), .input_share0(d3_P3_26_s0), .input_share1(d3_P3_26_s1), .output_share0(d4_P3_26_s0), .output_share1(d4_P3_26_s1));
  reg_module u_reg_P3_27_d4 (.clk(clk), .input_share0(d3_P3_27_s0), .input_share1(d3_P3_27_s1), .output_share0(d4_P3_27_s0), .output_share1(d4_P3_27_s1));
  reg_module u_reg_P3_28_d4 (.clk(clk), .input_share0(d3_P3_28_s0), .input_share1(d3_P3_28_s1), .output_share0(d4_P3_28_s0), .output_share1(d4_P3_28_s1));
  reg_module u_reg_P3_29_d4 (.clk(clk), .input_share0(d3_P3_29_s0), .input_share1(d3_P3_29_s1), .output_share0(d4_P3_29_s0), .output_share1(d4_P3_29_s1));
  reg_module u_reg_P3_30_d4 (.clk(clk), .input_share0(d3_P3_30_s0), .input_share1(d3_P3_30_s1), .output_share0(d4_P3_30_s0), .output_share1(d4_P3_30_s1));
  reg_module u_reg_P3_31_d4 (.clk(clk), .input_share0(d3_P3_31_s0), .input_share1(d3_P3_31_s1), .output_share0(d4_P3_31_s0), .output_share1(d4_P3_31_s1));
  xor_module u_xor_G3_10_d4 (.x_share0(d4_t67_s0), .x_share1(d4_t67_s1), .y_share0(d4_G2_10_s0), .y_share1(d4_G2_10_s1), .z_share0(d4_G3_10_s0), .z_share1(d4_G3_10_s1));
  xor_module u_xor_G3_11_d4 (.x_share0(d4_t68_s0), .x_share1(d4_t68_s1), .y_share0(d4_G2_11_s0), .y_share1(d4_G2_11_s1), .z_share0(d4_G3_11_s0), .z_share1(d4_G3_11_s1));
  xor_module u_xor_G3_12_d4 (.x_share0(d4_t69_s0), .x_share1(d4_t69_s1), .y_share0(d4_G2_12_s0), .y_share1(d4_G2_12_s1), .z_share0(d4_G3_12_s0), .z_share1(d4_G3_12_s1));
  xor_module u_xor_G3_13_d4 (.x_share0(d4_t70_s0), .x_share1(d4_t70_s1), .y_share0(d4_G2_13_s0), .y_share1(d4_G2_13_s1), .z_share0(d4_G3_13_s0), .z_share1(d4_G3_13_s1));
  xor_module u_xor_G3_14_d4 (.x_share0(d4_t71_s0), .x_share1(d4_t71_s1), .y_share0(d4_G2_14_s0), .y_share1(d4_G2_14_s1), .z_share0(d4_G3_14_s0), .z_share1(d4_G3_14_s1));
  xor_module u_xor_G3_15_d4 (.x_share0(d4_t72_s0), .x_share1(d4_t72_s1), .y_share0(d4_G2_15_s0), .y_share1(d4_G2_15_s1), .z_share0(d4_G3_15_s0), .z_share1(d4_G3_15_s1));
  xor_module u_xor_G3_16_d4 (.x_share0(d4_t73_s0), .x_share1(d4_t73_s1), .y_share0(d4_G2_16_s0), .y_share1(d4_G2_16_s1), .z_share0(d4_G3_16_s0), .z_share1(d4_G3_16_s1));
  xor_module u_xor_G3_17_d4 (.x_share0(d4_t74_s0), .x_share1(d4_t74_s1), .y_share0(d4_G2_17_s0), .y_share1(d4_G2_17_s1), .z_share0(d4_G3_17_s0), .z_share1(d4_G3_17_s1));
  xor_module u_xor_G3_18_d4 (.x_share0(d4_t75_s0), .x_share1(d4_t75_s1), .y_share0(d4_G2_18_s0), .y_share1(d4_G2_18_s1), .z_share0(d4_G3_18_s0), .z_share1(d4_G3_18_s1));
  xor_module u_xor_G3_19_d4 (.x_share0(d4_t76_s0), .x_share1(d4_t76_s1), .y_share0(d4_G2_19_s0), .y_share1(d4_G2_19_s1), .z_share0(d4_G3_19_s0), .z_share1(d4_G3_19_s1));
  xor_module u_xor_G3_20_d4 (.x_share0(d4_t77_s0), .x_share1(d4_t77_s1), .y_share0(d4_G2_20_s0), .y_share1(d4_G2_20_s1), .z_share0(d4_G3_20_s0), .z_share1(d4_G3_20_s1));
  xor_module u_xor_G3_21_d4 (.x_share0(d4_t78_s0), .x_share1(d4_t78_s1), .y_share0(d4_G2_21_s0), .y_share1(d4_G2_21_s1), .z_share0(d4_G3_21_s0), .z_share1(d4_G3_21_s1));
  xor_module u_xor_G3_22_d4 (.x_share0(d4_t79_s0), .x_share1(d4_t79_s1), .y_share0(d4_G2_22_s0), .y_share1(d4_G2_22_s1), .z_share0(d4_G3_22_s0), .z_share1(d4_G3_22_s1));
  xor_module u_xor_G3_23_d4 (.x_share0(d4_t80_s0), .x_share1(d4_t80_s1), .y_share0(d4_G2_23_s0), .y_share1(d4_G2_23_s1), .z_share0(d4_G3_23_s0), .z_share1(d4_G3_23_s1));
  xor_module u_xor_G3_24_d4 (.x_share0(d4_t81_s0), .x_share1(d4_t81_s1), .y_share0(d4_G2_24_s0), .y_share1(d4_G2_24_s1), .z_share0(d4_G3_24_s0), .z_share1(d4_G3_24_s1));
  xor_module u_xor_G3_25_d4 (.x_share0(d4_t82_s0), .x_share1(d4_t82_s1), .y_share0(d4_G2_25_s0), .y_share1(d4_G2_25_s1), .z_share0(d4_G3_25_s0), .z_share1(d4_G3_25_s1));
  xor_module u_xor_G3_26_d4 (.x_share0(d4_t83_s0), .x_share1(d4_t83_s1), .y_share0(d4_G2_26_s0), .y_share1(d4_G2_26_s1), .z_share0(d4_G3_26_s0), .z_share1(d4_G3_26_s1));
  xor_module u_xor_G3_27_d4 (.x_share0(d4_t84_s0), .x_share1(d4_t84_s1), .y_share0(d4_G2_27_s0), .y_share1(d4_G2_27_s1), .z_share0(d4_G3_27_s0), .z_share1(d4_G3_27_s1));
  xor_module u_xor_G3_28_d4 (.x_share0(d4_t85_s0), .x_share1(d4_t85_s1), .y_share0(d4_G2_28_s0), .y_share1(d4_G2_28_s1), .z_share0(d4_G3_28_s0), .z_share1(d4_G3_28_s1));
  xor_module u_xor_G3_29_d4 (.x_share0(d4_t86_s0), .x_share1(d4_t86_s1), .y_share0(d4_G2_29_s0), .y_share1(d4_G2_29_s1), .z_share0(d4_G3_29_s0), .z_share1(d4_G3_29_s1));
  xor_module u_xor_G3_30_d4 (.x_share0(d4_t87_s0), .x_share1(d4_t87_s1), .y_share0(d4_G2_30_s0), .y_share1(d4_G2_30_s1), .z_share0(d4_G3_30_s0), .z_share1(d4_G3_30_s1));
  xor_module u_xor_G3_31_d4 (.x_share0(d4_t88_s0), .x_share1(d4_t88_s1), .y_share0(d4_G2_31_s0), .y_share1(d4_G2_31_s1), .z_share0(d4_G3_31_s0), .z_share1(d4_G3_31_s1));
  xor_module u_xor_G3_7_d4 (.x_share0(d4_t64_s0), .x_share1(d4_t64_s1), .y_share0(d4_G2_7_s0), .y_share1(d4_G2_7_s1), .z_share0(d4_G3_7_s0), .z_share1(d4_G3_7_s1));
  xor_module u_xor_G3_8_d4 (.x_share0(d4_t65_s0), .x_share1(d4_t65_s1), .y_share0(d4_G2_8_s0), .y_share1(d4_G2_8_s1), .z_share0(d4_G3_8_s0), .z_share1(d4_G3_8_s1));
  xor_module u_xor_G3_9_d4 (.x_share0(d4_t66_s0), .x_share1(d4_t66_s1), .y_share0(d4_G2_9_s0), .y_share1(d4_G2_9_s1), .z_share0(d4_G3_9_s0), .z_share1(d4_G3_9_s1));
  xor_module u_xor_G4_10_d4 (.x_share0(d4_t91_s0), .x_share1(d4_t91_s1), .y_share0(d4_G3_10_s0), .y_share1(d4_G3_10_s1), .z_share0(d4_G4_10_s0), .z_share1(d4_G4_10_s1));
  xor_module u_xor_G4_11_d4 (.x_share0(d4_t92_s0), .x_share1(d4_t92_s1), .y_share0(d4_G3_11_s0), .y_share1(d4_G3_11_s1), .z_share0(d4_G4_11_s0), .z_share1(d4_G4_11_s1));
  xor_module u_xor_G4_12_d4 (.x_share0(d4_t93_s0), .x_share1(d4_t93_s1), .y_share0(d4_G3_12_s0), .y_share1(d4_G3_12_s1), .z_share0(d4_G4_12_s0), .z_share1(d4_G4_12_s1));
  xor_module u_xor_G4_13_d4 (.x_share0(d4_t94_s0), .x_share1(d4_t94_s1), .y_share0(d4_G3_13_s0), .y_share1(d4_G3_13_s1), .z_share0(d4_G4_13_s0), .z_share1(d4_G4_13_s1));
  xor_module u_xor_G4_14_d4 (.x_share0(d4_t95_s0), .x_share1(d4_t95_s1), .y_share0(d4_G3_14_s0), .y_share1(d4_G3_14_s1), .z_share0(d4_G4_14_s0), .z_share1(d4_G4_14_s1));
  xor_module u_xor_G4_8_d4 (.x_share0(d4_t89_s0), .x_share1(d4_t89_s1), .y_share0(d4_G3_8_s0), .y_share1(d4_G3_8_s1), .z_share0(d4_G4_8_s0), .z_share1(d4_G4_8_s1));
  xor_module u_xor_G4_9_d4 (.x_share0(d4_t90_s0), .x_share1(d4_t90_s1), .y_share0(d4_G3_9_s0), .y_share1(d4_G3_9_s1), .z_share0(d4_G4_9_s0), .z_share1(d4_G4_9_s1));
  and_module u_and_P4_16_d4 (.clk(clk), .x_share0(d3_P3_16_s0), .x_share1(d3_P3_16_s1), .y_share0(d3_P3_8_s0), .y_share1(d3_P3_8_s1), .rand(r_P4_16), .z_share0(d4_P4_16_s0), .z_share1(d4_P4_16_s1));
  assign r_P4_16 = stage4_share0[8];
  and_module u_and_P4_17_d4 (.clk(clk), .x_share0(d3_P3_17_s0), .x_share1(d3_P3_17_s1), .y_share0(d3_P3_9_s0), .y_share1(d3_P3_9_s1), .rand(r_P4_17), .z_share0(d4_P4_17_s0), .z_share1(d4_P4_17_s1));
  assign r_P4_17 = stage4_share0[4];
  and_module u_and_P4_18_d4 (.clk(clk), .x_share0(d3_P3_18_s0), .x_share1(d3_P3_18_s1), .y_share0(d3_P3_10_s0), .y_share1(d3_P3_10_s1), .rand(r_P4_18), .z_share0(d4_P4_18_s0), .z_share1(d4_P4_18_s1));
  assign r_P4_18 = stage4_share0[15];
  and_module u_and_P4_19_d4 (.clk(clk), .x_share0(d3_P3_19_s0), .x_share1(d3_P3_19_s1), .y_share0(d3_P3_11_s0), .y_share1(d3_P3_11_s1), .rand(r_P4_19), .z_share0(d4_P4_19_s0), .z_share1(d4_P4_19_s1));
  assign r_P4_19 = stage4_share0[9];
  and_module u_and_P4_20_d4 (.clk(clk), .x_share0(d3_P3_20_s0), .x_share1(d3_P3_20_s1), .y_share0(d3_P3_12_s0), .y_share1(d3_P3_12_s1), .rand(r_P4_20), .z_share0(d4_P4_20_s0), .z_share1(d4_P4_20_s1));
  assign r_P4_20 = stage4_share0[8];
  and_module u_and_P4_21_d4 (.clk(clk), .x_share0(d3_P3_21_s0), .x_share1(d3_P3_21_s1), .y_share0(d3_P3_13_s0), .y_share1(d3_P3_13_s1), .rand(r_P4_21), .z_share0(d4_P4_21_s0), .z_share1(d4_P4_21_s1));
  assign r_P4_21 = stage4_share0[4];
  and_module u_and_P4_22_d4 (.clk(clk), .x_share0(d3_P3_22_s0), .x_share1(d3_P3_22_s1), .y_share0(d3_P3_14_s0), .y_share1(d3_P3_14_s1), .rand(r_P4_22), .z_share0(d4_P4_22_s0), .z_share1(d4_P4_22_s1));
  assign r_P4_22 = stage4_share0[18];
  and_module u_and_P4_23_d4 (.clk(clk), .x_share0(d3_P3_23_s0), .x_share1(d3_P3_23_s1), .y_share0(d3_P3_15_s0), .y_share1(d3_P3_15_s1), .rand(r_P4_23), .z_share0(d4_P4_23_s0), .z_share1(d4_P4_23_s1));
  assign r_P4_23 = stage4_share0[9];
  and_module u_and_P4_24_d4 (.clk(clk), .x_share0(d3_P3_24_s0), .x_share1(d3_P3_24_s1), .y_share0(d3_P3_16_s0), .y_share1(d3_P3_16_s1), .rand(r_P4_24), .z_share0(d4_P4_24_s0), .z_share1(d4_P4_24_s1));
  assign r_P4_24 = stage4_share0[19];
  and_module u_and_P4_25_d4 (.clk(clk), .x_share0(d3_P3_25_s0), .x_share1(d3_P3_25_s1), .y_share0(d3_P3_17_s0), .y_share1(d3_P3_17_s1), .rand(r_P4_25), .z_share0(d4_P4_25_s0), .z_share1(d4_P4_25_s1));
  assign r_P4_25 = stage4_share0[21];
  and_module u_and_P4_26_d4 (.clk(clk), .x_share0(d3_P3_26_s0), .x_share1(d3_P3_26_s1), .y_share0(d3_P3_18_s0), .y_share1(d3_P3_18_s1), .rand(r_P4_26), .z_share0(d4_P4_26_s0), .z_share1(d4_P4_26_s1));
  assign r_P4_26 = stage4_share0[19];
  and_module u_and_P4_27_d4 (.clk(clk), .x_share0(d3_P3_27_s0), .x_share1(d3_P3_27_s1), .y_share0(d3_P3_19_s0), .y_share1(d3_P3_19_s1), .rand(r_P4_27), .z_share0(d4_P4_27_s0), .z_share1(d4_P4_27_s1));
  assign r_P4_27 = stage4_share0[23];
  and_module u_and_P4_28_d4 (.clk(clk), .x_share0(d3_P3_28_s0), .x_share1(d3_P3_28_s1), .y_share0(d3_P3_20_s0), .y_share1(d3_P3_20_s1), .rand(r_P4_28), .z_share0(d4_P4_28_s0), .z_share1(d4_P4_28_s1));
  assign r_P4_28 = stage4_share0[22];
  and_module u_and_P4_29_d4 (.clk(clk), .x_share0(d3_P3_29_s0), .x_share1(d3_P3_29_s1), .y_share0(d3_P3_21_s0), .y_share1(d3_P3_21_s1), .rand(r_P4_29), .z_share0(d4_P4_29_s0), .z_share1(d4_P4_29_s1));
  assign r_P4_29 = stage4_share0[24];
  and_module u_and_P4_30_d4 (.clk(clk), .x_share0(d3_P3_30_s0), .x_share1(d3_P3_30_s1), .y_share0(d3_P3_22_s0), .y_share1(d3_P3_22_s1), .rand(r_P4_30), .z_share0(d4_P4_30_s0), .z_share1(d4_P4_30_s1));
  assign r_P4_30 = stage4_share0[24];
  and_module u_and_P4_31_d4 (.clk(clk), .x_share0(d3_P3_31_s0), .x_share1(d3_P3_31_s1), .y_share0(d3_P3_23_s0), .y_share1(d3_P3_23_s1), .rand(r_P4_31), .z_share0(d4_P4_31_s0), .z_share1(d4_P4_31_s1));
  assign r_P4_31 = stage4_share0[7];
  xor_module u_xor_o10_d4 (.x_share0(d4_P0_10_s0), .x_share1(d4_P0_10_s1), .y_share0(d4_G4_9_s0), .y_share1(d4_G4_9_s1), .z_share0(d4_o10_s0), .z_share1(d4_o10_s1));
  xor_module u_xor_o11_d4 (.x_share0(d4_P0_11_s0), .x_share1(d4_P0_11_s1), .y_share0(d4_G4_10_s0), .y_share1(d4_G4_10_s1), .z_share0(d4_o11_s0), .z_share1(d4_o11_s1));
  xor_module u_xor_o12_d4 (.x_share0(d4_P0_12_s0), .x_share1(d4_P0_12_s1), .y_share0(d4_G4_11_s0), .y_share1(d4_G4_11_s1), .z_share0(d4_o12_s0), .z_share1(d4_o12_s1));
  xor_module u_xor_o13_d4 (.x_share0(d4_P0_13_s0), .x_share1(d4_P0_13_s1), .y_share0(d4_G4_12_s0), .y_share1(d4_G4_12_s1), .z_share0(d4_o13_s0), .z_share1(d4_o13_s1));
  xor_module u_xor_o14_d4 (.x_share0(d4_P0_14_s0), .x_share1(d4_P0_14_s1), .y_share0(d4_G4_13_s0), .y_share1(d4_G4_13_s1), .z_share0(d4_o14_s0), .z_share1(d4_o14_s1));
  xor_module u_xor_o15_d4 (.x_share0(d4_P0_15_s0), .x_share1(d4_P0_15_s1), .y_share0(d4_G4_14_s0), .y_share1(d4_G4_14_s1), .z_share0(d4_o15_s0), .z_share1(d4_o15_s1));
  xor_module u_xor_o8_d4 (.x_share0(d4_P0_8_s0), .x_share1(d4_P0_8_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .z_share0(d4_o8_s0), .z_share1(d4_o8_s1));
  xor_module u_xor_o9_d4 (.x_share0(d4_P0_9_s0), .x_share1(d4_P0_9_s1), .y_share0(d4_G4_8_s0), .y_share1(d4_G4_8_s1), .z_share0(d4_o9_s0), .z_share1(d4_o9_s1));
  and_module u_and_t64_d4 (.clk(clk), .x_share0(d3_P2_7_s0), .x_share1(d3_P2_7_s1), .y_share0(d3_G2_3_s0), .y_share1(d3_G2_3_s1), .rand(r_t64), .z_share0(d4_t64_s0), .z_share1(d4_t64_s1));
  assign r_t64 = stage4_share0[22];
  and_module u_and_t65_d4 (.clk(clk), .x_share0(d3_P2_8_s0), .x_share1(d3_P2_8_s1), .y_share0(d3_G2_4_s0), .y_share1(d3_G2_4_s1), .rand(r_t65), .z_share0(d4_t65_s0), .z_share1(d4_t65_s1));
  assign r_t65 = stage4_share0[13];
  and_module u_and_t66_d4 (.clk(clk), .x_share0(d3_P2_9_s0), .x_share1(d3_P2_9_s1), .y_share0(d3_G2_5_s0), .y_share1(d3_G2_5_s1), .rand(r_t66), .z_share0(d4_t66_s0), .z_share1(d4_t66_s1));
  assign r_t66 = stage4_share0[15];
  and_module u_and_t67_d4 (.clk(clk), .x_share0(d3_P2_10_s0), .x_share1(d3_P2_10_s1), .y_share0(d3_G2_6_s0), .y_share1(d3_G2_6_s1), .rand(r_t67), .z_share0(d4_t67_s0), .z_share1(d4_t67_s1));
  assign r_t67 = stage4_share0[0];
  and_module u_and_t68_d4 (.clk(clk), .x_share0(d3_P2_11_s0), .x_share1(d3_P2_11_s1), .y_share0(d3_G2_7_s0), .y_share1(d3_G2_7_s1), .rand(r_t68), .z_share0(d4_t68_s0), .z_share1(d4_t68_s1));
  assign r_t68 = stage4_share0[8];
  and_module u_and_t69_d4 (.clk(clk), .x_share0(d3_P2_12_s0), .x_share1(d3_P2_12_s1), .y_share0(d3_G2_8_s0), .y_share1(d3_G2_8_s1), .rand(r_t69), .z_share0(d4_t69_s0), .z_share1(d4_t69_s1));
  assign r_t69 = stage4_share0[23];
  and_module u_and_t70_d4 (.clk(clk), .x_share0(d3_P2_13_s0), .x_share1(d3_P2_13_s1), .y_share0(d3_G2_9_s0), .y_share1(d3_G2_9_s1), .rand(r_t70), .z_share0(d4_t70_s0), .z_share1(d4_t70_s1));
  assign r_t70 = stage4_share0[3];
  and_module u_and_t71_d4 (.clk(clk), .x_share0(d3_P2_14_s0), .x_share1(d3_P2_14_s1), .y_share0(d3_G2_10_s0), .y_share1(d3_G2_10_s1), .rand(r_t71), .z_share0(d4_t71_s0), .z_share1(d4_t71_s1));
  assign r_t71 = stage4_share0[15];
  and_module u_and_t72_d4 (.clk(clk), .x_share0(d3_P2_15_s0), .x_share1(d3_P2_15_s1), .y_share0(d3_G2_11_s0), .y_share1(d3_G2_11_s1), .rand(r_t72), .z_share0(d4_t72_s0), .z_share1(d4_t72_s1));
  assign r_t72 = stage4_share0[5];
  and_module u_and_t73_d4 (.clk(clk), .x_share0(d3_P2_16_s0), .x_share1(d3_P2_16_s1), .y_share0(d3_G2_12_s0), .y_share1(d3_G2_12_s1), .rand(r_t73), .z_share0(d4_t73_s0), .z_share1(d4_t73_s1));
  assign r_t73 = stage4_share0[7];
  and_module u_and_t74_d4 (.clk(clk), .x_share0(d3_P2_17_s0), .x_share1(d3_P2_17_s1), .y_share0(d3_G2_13_s0), .y_share1(d3_G2_13_s1), .rand(r_t74), .z_share0(d4_t74_s0), .z_share1(d4_t74_s1));
  assign r_t74 = stage4_share0[19];
  and_module u_and_t75_d4 (.clk(clk), .x_share0(d3_P2_18_s0), .x_share1(d3_P2_18_s1), .y_share0(d3_G2_14_s0), .y_share1(d3_G2_14_s1), .rand(r_t75), .z_share0(d4_t75_s0), .z_share1(d4_t75_s1));
  assign r_t75 = stage4_share0[16];
  and_module u_and_t76_d4 (.clk(clk), .x_share0(d3_P2_19_s0), .x_share1(d3_P2_19_s1), .y_share0(d3_G2_15_s0), .y_share1(d3_G2_15_s1), .rand(r_t76), .z_share0(d4_t76_s0), .z_share1(d4_t76_s1));
  assign r_t76 = stage4_share0[19];
  and_module u_and_t77_d4 (.clk(clk), .x_share0(d3_P2_20_s0), .x_share1(d3_P2_20_s1), .y_share0(d3_G2_16_s0), .y_share1(d3_G2_16_s1), .rand(r_t77), .z_share0(d4_t77_s0), .z_share1(d4_t77_s1));
  assign r_t77 = stage4_share0[11];
  and_module u_and_t78_d4 (.clk(clk), .x_share0(d3_P2_21_s0), .x_share1(d3_P2_21_s1), .y_share0(d3_G2_17_s0), .y_share1(d3_G2_17_s1), .rand(r_t78), .z_share0(d4_t78_s0), .z_share1(d4_t78_s1));
  assign r_t78 = stage4_share0[10];
  and_module u_and_t79_d4 (.clk(clk), .x_share0(d3_P2_22_s0), .x_share1(d3_P2_22_s1), .y_share0(d3_G2_18_s0), .y_share1(d3_G2_18_s1), .rand(r_t79), .z_share0(d4_t79_s0), .z_share1(d4_t79_s1));
  assign r_t79 = stage4_share0[14];
  and_module u_and_t80_d4 (.clk(clk), .x_share0(d3_P2_23_s0), .x_share1(d3_P2_23_s1), .y_share0(d3_G2_19_s0), .y_share1(d3_G2_19_s1), .rand(r_t80), .z_share0(d4_t80_s0), .z_share1(d4_t80_s1));
  assign r_t80 = stage4_share0[10];
  and_module u_and_t81_d4 (.clk(clk), .x_share0(d3_P2_24_s0), .x_share1(d3_P2_24_s1), .y_share0(d3_G2_20_s0), .y_share1(d3_G2_20_s1), .rand(r_t81), .z_share0(d4_t81_s0), .z_share1(d4_t81_s1));
  assign r_t81 = stage4_share0[22];
  and_module u_and_t82_d4 (.clk(clk), .x_share0(d3_P2_25_s0), .x_share1(d3_P2_25_s1), .y_share0(d3_G2_21_s0), .y_share1(d3_G2_21_s1), .rand(r_t82), .z_share0(d4_t82_s0), .z_share1(d4_t82_s1));
  assign r_t82 = stage4_share0[23];
  and_module u_and_t83_d4 (.clk(clk), .x_share0(d3_P2_26_s0), .x_share1(d3_P2_26_s1), .y_share0(d3_G2_22_s0), .y_share1(d3_G2_22_s1), .rand(r_t83), .z_share0(d4_t83_s0), .z_share1(d4_t83_s1));
  assign r_t83 = stage4_share0[21];
  and_module u_and_t84_d4 (.clk(clk), .x_share0(d3_P2_27_s0), .x_share1(d3_P2_27_s1), .y_share0(d3_G2_23_s0), .y_share1(d3_G2_23_s1), .rand(r_t84), .z_share0(d4_t84_s0), .z_share1(d4_t84_s1));
  assign r_t84 = stage4_share0[22];
  and_module u_and_t85_d4 (.clk(clk), .x_share0(d3_P2_28_s0), .x_share1(d3_P2_28_s1), .y_share0(d3_G2_24_s0), .y_share1(d3_G2_24_s1), .rand(r_t85), .z_share0(d4_t85_s0), .z_share1(d4_t85_s1));
  assign r_t85 = stage4_share0[6];
  and_module u_and_t86_d4 (.clk(clk), .x_share0(d3_P2_29_s0), .x_share1(d3_P2_29_s1), .y_share0(d3_G2_25_s0), .y_share1(d3_G2_25_s1), .rand(r_t86), .z_share0(d4_t86_s0), .z_share1(d4_t86_s1));
  assign r_t86 = stage4_share0[14];
  and_module u_and_t87_d4 (.clk(clk), .x_share0(d3_P2_30_s0), .x_share1(d3_P2_30_s1), .y_share0(d3_G2_26_s0), .y_share1(d3_G2_26_s1), .rand(r_t87), .z_share0(d4_t87_s0), .z_share1(d4_t87_s1));
  assign r_t87 = stage4_share0[13];
  and_module u_and_t88_d4 (.clk(clk), .x_share0(d3_P2_31_s0), .x_share1(d3_P2_31_s1), .y_share0(d3_G2_27_s0), .y_share1(d3_G2_27_s1), .rand(r_t88), .z_share0(d4_t88_s0), .z_share1(d4_t88_s1));
  assign r_t88 = stage4_share0[12];
  and_module u_and_t89_d4 (.clk(clk), .x_share0(d3_P3_8_s0), .x_share1(d3_P3_8_s1), .y_share0(d3_G0_0_s0), .y_share1(d3_G0_0_s1), .rand(r_t89), .z_share0(d4_t89_s0), .z_share1(d4_t89_s1));
  assign r_t89 = stage4_share0[20];
  and_module u_and_t90_d4 (.clk(clk), .x_share0(d3_P3_9_s0), .x_share1(d3_P3_9_s1), .y_share0(d3_G1_1_s0), .y_share1(d3_G1_1_s1), .rand(r_t90), .z_share0(d4_t90_s0), .z_share1(d4_t90_s1));
  assign r_t90 = stage4_share0[17];
  and_module u_and_t91_d4 (.clk(clk), .x_share0(d3_P3_10_s0), .x_share1(d3_P3_10_s1), .y_share0(d3_G2_2_s0), .y_share1(d3_G2_2_s1), .rand(r_t91), .z_share0(d4_t91_s0), .z_share1(d4_t91_s1));
  assign r_t91 = stage4_share0[7];
  and_module u_and_t92_d4 (.clk(clk), .x_share0(d3_P3_11_s0), .x_share1(d3_P3_11_s1), .y_share0(d3_G2_3_s0), .y_share1(d3_G2_3_s1), .rand(r_t92), .z_share0(d4_t92_s0), .z_share1(d4_t92_s1));
  assign r_t92 = stage4_share0[11];
  and_module u_and_t93_d4 (.clk(clk), .x_share0(d3_P3_12_s0), .x_share1(d3_P3_12_s1), .y_share0(d3_G3_4_s0), .y_share1(d3_G3_4_s1), .rand(r_t93), .z_share0(d4_t93_s0), .z_share1(d4_t93_s1));
  assign r_t93 = stage4_share0[5];
  and_module u_and_t94_d4 (.clk(clk), .x_share0(d3_P3_13_s0), .x_share1(d3_P3_13_s1), .y_share0(d3_G3_5_s0), .y_share1(d3_G3_5_s1), .rand(r_t94), .z_share0(d4_t94_s0), .z_share1(d4_t94_s1));
  assign r_t94 = stage4_share0[25];
  and_module u_and_t95_d4 (.clk(clk), .x_share0(d3_P3_14_s0), .x_share1(d3_P3_14_s1), .y_share0(d3_G3_6_s0), .y_share1(d3_G3_6_s1), .rand(r_t95), .z_share0(d4_t95_s0), .z_share1(d4_t95_s1));
  assign r_t95 = stage4_share0[8];
  reg_module u_reg_G3_15_d5 (.clk(clk), .input_share0(d4_G3_15_s0), .input_share1(d4_G3_15_s1), .output_share0(d5_G3_15_s0), .output_share1(d5_G3_15_s1));
  reg_module u_reg_G3_16_d5 (.clk(clk), .input_share0(d4_G3_16_s0), .input_share1(d4_G3_16_s1), .output_share0(d5_G3_16_s0), .output_share1(d5_G3_16_s1));
  reg_module u_reg_G3_17_d5 (.clk(clk), .input_share0(d4_G3_17_s0), .input_share1(d4_G3_17_s1), .output_share0(d5_G3_17_s0), .output_share1(d5_G3_17_s1));
  reg_module u_reg_G3_18_d5 (.clk(clk), .input_share0(d4_G3_18_s0), .input_share1(d4_G3_18_s1), .output_share0(d5_G3_18_s0), .output_share1(d5_G3_18_s1));
  reg_module u_reg_G3_19_d5 (.clk(clk), .input_share0(d4_G3_19_s0), .input_share1(d4_G3_19_s1), .output_share0(d5_G3_19_s0), .output_share1(d5_G3_19_s1));
  reg_module u_reg_G3_20_d5 (.clk(clk), .input_share0(d4_G3_20_s0), .input_share1(d4_G3_20_s1), .output_share0(d5_G3_20_s0), .output_share1(d5_G3_20_s1));
  reg_module u_reg_G3_21_d5 (.clk(clk), .input_share0(d4_G3_21_s0), .input_share1(d4_G3_21_s1), .output_share0(d5_G3_21_s0), .output_share1(d5_G3_21_s1));
  reg_module u_reg_G3_22_d5 (.clk(clk), .input_share0(d4_G3_22_s0), .input_share1(d4_G3_22_s1), .output_share0(d5_G3_22_s0), .output_share1(d5_G3_22_s1));
  reg_module u_reg_G3_23_d5 (.clk(clk), .input_share0(d4_G3_23_s0), .input_share1(d4_G3_23_s1), .output_share0(d5_G3_23_s0), .output_share1(d5_G3_23_s1));
  reg_module u_reg_G3_24_d5 (.clk(clk), .input_share0(d4_G3_24_s0), .input_share1(d4_G3_24_s1), .output_share0(d5_G3_24_s0), .output_share1(d5_G3_24_s1));
  reg_module u_reg_G3_25_d5 (.clk(clk), .input_share0(d4_G3_25_s0), .input_share1(d4_G3_25_s1), .output_share0(d5_G3_25_s0), .output_share1(d5_G3_25_s1));
  reg_module u_reg_G3_26_d5 (.clk(clk), .input_share0(d4_G3_26_s0), .input_share1(d4_G3_26_s1), .output_share0(d5_G3_26_s0), .output_share1(d5_G3_26_s1));
  reg_module u_reg_G3_27_d5 (.clk(clk), .input_share0(d4_G3_27_s0), .input_share1(d4_G3_27_s1), .output_share0(d5_G3_27_s0), .output_share1(d5_G3_27_s1));
  reg_module u_reg_G3_28_d5 (.clk(clk), .input_share0(d4_G3_28_s0), .input_share1(d4_G3_28_s1), .output_share0(d5_G3_28_s0), .output_share1(d5_G3_28_s1));
  reg_module u_reg_G3_29_d5 (.clk(clk), .input_share0(d4_G3_29_s0), .input_share1(d4_G3_29_s1), .output_share0(d5_G3_29_s0), .output_share1(d5_G3_29_s1));
  reg_module u_reg_G3_30_d5 (.clk(clk), .input_share0(d4_G3_30_s0), .input_share1(d4_G3_30_s1), .output_share0(d5_G3_30_s0), .output_share1(d5_G3_30_s1));
  reg_module u_reg_G3_31_d5 (.clk(clk), .input_share0(d4_G3_31_s0), .input_share1(d4_G3_31_s1), .output_share0(d5_G3_31_s0), .output_share1(d5_G3_31_s1));
  reg_module u_reg_P0_16_d5 (.clk(clk), .input_share0(d4_P0_16_s0), .input_share1(d4_P0_16_s1), .output_share0(d5_P0_16_s0), .output_share1(d5_P0_16_s1));
  reg_module u_reg_P0_17_d5 (.clk(clk), .input_share0(d4_P0_17_s0), .input_share1(d4_P0_17_s1), .output_share0(d5_P0_17_s0), .output_share1(d5_P0_17_s1));
  reg_module u_reg_P0_18_d5 (.clk(clk), .input_share0(d4_P0_18_s0), .input_share1(d4_P0_18_s1), .output_share0(d5_P0_18_s0), .output_share1(d5_P0_18_s1));
  reg_module u_reg_P0_19_d5 (.clk(clk), .input_share0(d4_P0_19_s0), .input_share1(d4_P0_19_s1), .output_share0(d5_P0_19_s0), .output_share1(d5_P0_19_s1));
  reg_module u_reg_P0_20_d5 (.clk(clk), .input_share0(d4_P0_20_s0), .input_share1(d4_P0_20_s1), .output_share0(d5_P0_20_s0), .output_share1(d5_P0_20_s1));
  reg_module u_reg_P0_21_d5 (.clk(clk), .input_share0(d4_P0_21_s0), .input_share1(d4_P0_21_s1), .output_share0(d5_P0_21_s0), .output_share1(d5_P0_21_s1));
  reg_module u_reg_P0_22_d5 (.clk(clk), .input_share0(d4_P0_22_s0), .input_share1(d4_P0_22_s1), .output_share0(d5_P0_22_s0), .output_share1(d5_P0_22_s1));
  reg_module u_reg_P0_23_d5 (.clk(clk), .input_share0(d4_P0_23_s0), .input_share1(d4_P0_23_s1), .output_share0(d5_P0_23_s0), .output_share1(d5_P0_23_s1));
  reg_module u_reg_P0_24_d5 (.clk(clk), .input_share0(d4_P0_24_s0), .input_share1(d4_P0_24_s1), .output_share0(d5_P0_24_s0), .output_share1(d5_P0_24_s1));
  reg_module u_reg_P0_25_d5 (.clk(clk), .input_share0(d4_P0_25_s0), .input_share1(d4_P0_25_s1), .output_share0(d5_P0_25_s0), .output_share1(d5_P0_25_s1));
  reg_module u_reg_P0_26_d5 (.clk(clk), .input_share0(d4_P0_26_s0), .input_share1(d4_P0_26_s1), .output_share0(d5_P0_26_s0), .output_share1(d5_P0_26_s1));
  reg_module u_reg_P0_27_d5 (.clk(clk), .input_share0(d4_P0_27_s0), .input_share1(d4_P0_27_s1), .output_share0(d5_P0_27_s0), .output_share1(d5_P0_27_s1));
  reg_module u_reg_P0_28_d5 (.clk(clk), .input_share0(d4_P0_28_s0), .input_share1(d4_P0_28_s1), .output_share0(d5_P0_28_s0), .output_share1(d5_P0_28_s1));
  reg_module u_reg_P0_29_d5 (.clk(clk), .input_share0(d4_P0_29_s0), .input_share1(d4_P0_29_s1), .output_share0(d5_P0_29_s0), .output_share1(d5_P0_29_s1));
  reg_module u_reg_P0_30_d5 (.clk(clk), .input_share0(d4_P0_30_s0), .input_share1(d4_P0_30_s1), .output_share0(d5_P0_30_s0), .output_share1(d5_P0_30_s1));
  reg_module u_reg_P0_31_d5 (.clk(clk), .input_share0(d4_P0_31_s0), .input_share1(d4_P0_31_s1), .output_share0(d5_P0_31_s0), .output_share1(d5_P0_31_s1));
  reg_module u_reg_P4_31_d5 (.clk(clk), .input_share0(d4_P4_31_s0), .input_share1(d4_P4_31_s1), .output_share0(d5_P4_31_s0), .output_share1(d5_P4_31_s1));
  xor_module u_xor_G4_15_d5 (.x_share0(d5_t96_s0), .x_share1(d5_t96_s1), .y_share0(d5_G3_15_s0), .y_share1(d5_G3_15_s1), .z_share0(d5_G4_15_s0), .z_share1(d5_G4_15_s1));
  xor_module u_xor_G4_16_d5 (.x_share0(d5_t97_s0), .x_share1(d5_t97_s1), .y_share0(d5_G3_16_s0), .y_share1(d5_G3_16_s1), .z_share0(d5_G4_16_s0), .z_share1(d5_G4_16_s1));
  xor_module u_xor_G4_17_d5 (.x_share0(d5_t98_s0), .x_share1(d5_t98_s1), .y_share0(d5_G3_17_s0), .y_share1(d5_G3_17_s1), .z_share0(d5_G4_17_s0), .z_share1(d5_G4_17_s1));
  xor_module u_xor_G4_18_d5 (.x_share0(d5_t99_s0), .x_share1(d5_t99_s1), .y_share0(d5_G3_18_s0), .y_share1(d5_G3_18_s1), .z_share0(d5_G4_18_s0), .z_share1(d5_G4_18_s1));
  xor_module u_xor_G4_19_d5 (.x_share0(d5_t100_s0), .x_share1(d5_t100_s1), .y_share0(d5_G3_19_s0), .y_share1(d5_G3_19_s1), .z_share0(d5_G4_19_s0), .z_share1(d5_G4_19_s1));
  xor_module u_xor_G4_20_d5 (.x_share0(d5_t101_s0), .x_share1(d5_t101_s1), .y_share0(d5_G3_20_s0), .y_share1(d5_G3_20_s1), .z_share0(d5_G4_20_s0), .z_share1(d5_G4_20_s1));
  xor_module u_xor_G4_21_d5 (.x_share0(d5_t102_s0), .x_share1(d5_t102_s1), .y_share0(d5_G3_21_s0), .y_share1(d5_G3_21_s1), .z_share0(d5_G4_21_s0), .z_share1(d5_G4_21_s1));
  xor_module u_xor_G4_22_d5 (.x_share0(d5_t103_s0), .x_share1(d5_t103_s1), .y_share0(d5_G3_22_s0), .y_share1(d5_G3_22_s1), .z_share0(d5_G4_22_s0), .z_share1(d5_G4_22_s1));
  xor_module u_xor_G4_23_d5 (.x_share0(d5_t104_s0), .x_share1(d5_t104_s1), .y_share0(d5_G3_23_s0), .y_share1(d5_G3_23_s1), .z_share0(d5_G4_23_s0), .z_share1(d5_G4_23_s1));
  xor_module u_xor_G4_24_d5 (.x_share0(d5_t105_s0), .x_share1(d5_t105_s1), .y_share0(d5_G3_24_s0), .y_share1(d5_G3_24_s1), .z_share0(d5_G4_24_s0), .z_share1(d5_G4_24_s1));
  xor_module u_xor_G4_25_d5 (.x_share0(d5_t106_s0), .x_share1(d5_t106_s1), .y_share0(d5_G3_25_s0), .y_share1(d5_G3_25_s1), .z_share0(d5_G4_25_s0), .z_share1(d5_G4_25_s1));
  xor_module u_xor_G4_26_d5 (.x_share0(d5_t107_s0), .x_share1(d5_t107_s1), .y_share0(d5_G3_26_s0), .y_share1(d5_G3_26_s1), .z_share0(d5_G4_26_s0), .z_share1(d5_G4_26_s1));
  xor_module u_xor_G4_27_d5 (.x_share0(d5_t108_s0), .x_share1(d5_t108_s1), .y_share0(d5_G3_27_s0), .y_share1(d5_G3_27_s1), .z_share0(d5_G4_27_s0), .z_share1(d5_G4_27_s1));
  xor_module u_xor_G4_28_d5 (.x_share0(d5_t109_s0), .x_share1(d5_t109_s1), .y_share0(d5_G3_28_s0), .y_share1(d5_G3_28_s1), .z_share0(d5_G4_28_s0), .z_share1(d5_G4_28_s1));
  xor_module u_xor_G4_29_d5 (.x_share0(d5_t110_s0), .x_share1(d5_t110_s1), .y_share0(d5_G3_29_s0), .y_share1(d5_G3_29_s1), .z_share0(d5_G4_29_s0), .z_share1(d5_G4_29_s1));
  xor_module u_xor_G4_30_d5 (.x_share0(d5_t111_s0), .x_share1(d5_t111_s1), .y_share0(d5_G3_30_s0), .y_share1(d5_G3_30_s1), .z_share0(d5_G4_30_s0), .z_share1(d5_G4_30_s1));
  xor_module u_xor_G4_31_d5 (.x_share0(d5_t112_s0), .x_share1(d5_t112_s1), .y_share0(d5_G3_31_s0), .y_share1(d5_G3_31_s1), .z_share0(d5_G4_31_s0), .z_share1(d5_G4_31_s1));
  xor_module u_xor_G5_16_d5 (.x_share0(d5_t113_s0), .x_share1(d5_t113_s1), .y_share0(d5_G4_16_s0), .y_share1(d5_G4_16_s1), .z_share0(d5_G5_16_s0), .z_share1(d5_G5_16_s1));
  xor_module u_xor_G5_17_d5 (.x_share0(d5_t114_s0), .x_share1(d5_t114_s1), .y_share0(d5_G4_17_s0), .y_share1(d5_G4_17_s1), .z_share0(d5_G5_17_s0), .z_share1(d5_G5_17_s1));
  xor_module u_xor_G5_18_d5 (.x_share0(d5_t115_s0), .x_share1(d5_t115_s1), .y_share0(d5_G4_18_s0), .y_share1(d5_G4_18_s1), .z_share0(d5_G5_18_s0), .z_share1(d5_G5_18_s1));
  xor_module u_xor_G5_19_d5 (.x_share0(d5_t116_s0), .x_share1(d5_t116_s1), .y_share0(d5_G4_19_s0), .y_share1(d5_G4_19_s1), .z_share0(d5_G5_19_s0), .z_share1(d5_G5_19_s1));
  xor_module u_xor_G5_20_d5 (.x_share0(d5_t117_s0), .x_share1(d5_t117_s1), .y_share0(d5_G4_20_s0), .y_share1(d5_G4_20_s1), .z_share0(d5_G5_20_s0), .z_share1(d5_G5_20_s1));
  xor_module u_xor_G5_21_d5 (.x_share0(d5_t118_s0), .x_share1(d5_t118_s1), .y_share0(d5_G4_21_s0), .y_share1(d5_G4_21_s1), .z_share0(d5_G5_21_s0), .z_share1(d5_G5_21_s1));
  xor_module u_xor_G5_22_d5 (.x_share0(d5_t119_s0), .x_share1(d5_t119_s1), .y_share0(d5_G4_22_s0), .y_share1(d5_G4_22_s1), .z_share0(d5_G5_22_s0), .z_share1(d5_G5_22_s1));
  xor_module u_xor_G5_23_d5 (.x_share0(d5_t120_s0), .x_share1(d5_t120_s1), .y_share0(d5_G4_23_s0), .y_share1(d5_G4_23_s1), .z_share0(d5_G5_23_s0), .z_share1(d5_G5_23_s1));
  xor_module u_xor_G5_24_d5 (.x_share0(d5_t121_s0), .x_share1(d5_t121_s1), .y_share0(d5_G4_24_s0), .y_share1(d5_G4_24_s1), .z_share0(d5_G5_24_s0), .z_share1(d5_G5_24_s1));
  xor_module u_xor_G5_25_d5 (.x_share0(d5_t122_s0), .x_share1(d5_t122_s1), .y_share0(d5_G4_25_s0), .y_share1(d5_G4_25_s1), .z_share0(d5_G5_25_s0), .z_share1(d5_G5_25_s1));
  xor_module u_xor_G5_26_d5 (.x_share0(d5_t123_s0), .x_share1(d5_t123_s1), .y_share0(d5_G4_26_s0), .y_share1(d5_G4_26_s1), .z_share0(d5_G5_26_s0), .z_share1(d5_G5_26_s1));
  xor_module u_xor_G5_27_d5 (.x_share0(d5_t124_s0), .x_share1(d5_t124_s1), .y_share0(d5_G4_27_s0), .y_share1(d5_G4_27_s1), .z_share0(d5_G5_27_s0), .z_share1(d5_G5_27_s1));
  xor_module u_xor_G5_28_d5 (.x_share0(d5_t125_s0), .x_share1(d5_t125_s1), .y_share0(d5_G4_28_s0), .y_share1(d5_G4_28_s1), .z_share0(d5_G5_28_s0), .z_share1(d5_G5_28_s1));
  xor_module u_xor_G5_29_d5 (.x_share0(d5_t126_s0), .x_share1(d5_t126_s1), .y_share0(d5_G4_29_s0), .y_share1(d5_G4_29_s1), .z_share0(d5_G5_29_s0), .z_share1(d5_G5_29_s1));
  xor_module u_xor_G5_30_d5 (.x_share0(d5_t127_s0), .x_share1(d5_t127_s1), .y_share0(d5_G4_30_s0), .y_share1(d5_G4_30_s1), .z_share0(d5_G5_30_s0), .z_share1(d5_G5_30_s1));
  xor_module u_xor_o16_d5 (.x_share0(d5_P0_16_s0), .x_share1(d5_P0_16_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .z_share0(d5_o16_s0), .z_share1(d5_o16_s1));
  xor_module u_xor_o17_d5 (.x_share0(d5_P0_17_s0), .x_share1(d5_P0_17_s1), .y_share0(d5_G5_16_s0), .y_share1(d5_G5_16_s1), .z_share0(d5_o17_s0), .z_share1(d5_o17_s1));
  xor_module u_xor_o18_d5 (.x_share0(d5_P0_18_s0), .x_share1(d5_P0_18_s1), .y_share0(d5_G5_17_s0), .y_share1(d5_G5_17_s1), .z_share0(d5_o18_s0), .z_share1(d5_o18_s1));
  xor_module u_xor_o19_d5 (.x_share0(d5_P0_19_s0), .x_share1(d5_P0_19_s1), .y_share0(d5_G5_18_s0), .y_share1(d5_G5_18_s1), .z_share0(d5_o19_s0), .z_share1(d5_o19_s1));
  xor_module u_xor_o20_d5 (.x_share0(d5_P0_20_s0), .x_share1(d5_P0_20_s1), .y_share0(d5_G5_19_s0), .y_share1(d5_G5_19_s1), .z_share0(d5_o20_s0), .z_share1(d5_o20_s1));
  xor_module u_xor_o21_d5 (.x_share0(d5_P0_21_s0), .x_share1(d5_P0_21_s1), .y_share0(d5_G5_20_s0), .y_share1(d5_G5_20_s1), .z_share0(d5_o21_s0), .z_share1(d5_o21_s1));
  xor_module u_xor_o22_d5 (.x_share0(d5_P0_22_s0), .x_share1(d5_P0_22_s1), .y_share0(d5_G5_21_s0), .y_share1(d5_G5_21_s1), .z_share0(d5_o22_s0), .z_share1(d5_o22_s1));
  xor_module u_xor_o23_d5 (.x_share0(d5_P0_23_s0), .x_share1(d5_P0_23_s1), .y_share0(d5_G5_22_s0), .y_share1(d5_G5_22_s1), .z_share0(d5_o23_s0), .z_share1(d5_o23_s1));
  xor_module u_xor_o24_d5 (.x_share0(d5_P0_24_s0), .x_share1(d5_P0_24_s1), .y_share0(d5_G5_23_s0), .y_share1(d5_G5_23_s1), .z_share0(d5_o24_s0), .z_share1(d5_o24_s1));
  xor_module u_xor_o25_d5 (.x_share0(d5_P0_25_s0), .x_share1(d5_P0_25_s1), .y_share0(d5_G5_24_s0), .y_share1(d5_G5_24_s1), .z_share0(d5_o25_s0), .z_share1(d5_o25_s1));
  xor_module u_xor_o26_d5 (.x_share0(d5_P0_26_s0), .x_share1(d5_P0_26_s1), .y_share0(d5_G5_25_s0), .y_share1(d5_G5_25_s1), .z_share0(d5_o26_s0), .z_share1(d5_o26_s1));
  xor_module u_xor_o27_d5 (.x_share0(d5_P0_27_s0), .x_share1(d5_P0_27_s1), .y_share0(d5_G5_26_s0), .y_share1(d5_G5_26_s1), .z_share0(d5_o27_s0), .z_share1(d5_o27_s1));
  xor_module u_xor_o28_d5 (.x_share0(d5_P0_28_s0), .x_share1(d5_P0_28_s1), .y_share0(d5_G5_27_s0), .y_share1(d5_G5_27_s1), .z_share0(d5_o28_s0), .z_share1(d5_o28_s1));
  xor_module u_xor_o29_d5 (.x_share0(d5_P0_29_s0), .x_share1(d5_P0_29_s1), .y_share0(d5_G5_28_s0), .y_share1(d5_G5_28_s1), .z_share0(d5_o29_s0), .z_share1(d5_o29_s1));
  xor_module u_xor_o30_d5 (.x_share0(d5_P0_30_s0), .x_share1(d5_P0_30_s1), .y_share0(d5_G5_29_s0), .y_share1(d5_G5_29_s1), .z_share0(d5_o30_s0), .z_share1(d5_o30_s1));
  xor_module u_xor_o31_d5 (.x_share0(d5_P0_31_s0), .x_share1(d5_P0_31_s1), .y_share0(d5_G5_30_s0), .y_share1(d5_G5_30_s1), .z_share0(d5_o31_s0), .z_share1(d5_o31_s1));
  and_module u_and_t100_d5 (.clk(clk), .x_share0(d4_P3_19_s0), .x_share1(d4_P3_19_s1), .y_share0(d4_G3_11_s0), .y_share1(d4_G3_11_s1), .rand(r_t100), .z_share0(d5_t100_s0), .z_share1(d5_t100_s1));
  assign r_t100 = stage5_share0[6];
  and_module u_and_t101_d5 (.clk(clk), .x_share0(d4_P3_20_s0), .x_share1(d4_P3_20_s1), .y_share0(d4_G3_12_s0), .y_share1(d4_G3_12_s1), .rand(r_t101), .z_share0(d5_t101_s0), .z_share1(d5_t101_s1));
  assign r_t101 = stage5_share0[18];
  and_module u_and_t102_d5 (.clk(clk), .x_share0(d4_P3_21_s0), .x_share1(d4_P3_21_s1), .y_share0(d4_G3_13_s0), .y_share1(d4_G3_13_s1), .rand(r_t102), .z_share0(d5_t102_s0), .z_share1(d5_t102_s1));
  assign r_t102 = stage5_share0[18];
  and_module u_and_t103_d5 (.clk(clk), .x_share0(d4_P3_22_s0), .x_share1(d4_P3_22_s1), .y_share0(d4_G3_14_s0), .y_share1(d4_G3_14_s1), .rand(r_t103), .z_share0(d5_t103_s0), .z_share1(d5_t103_s1));
  assign r_t103 = stage5_share0[9];
  and_module u_and_t104_d5 (.clk(clk), .x_share0(d4_P3_23_s0), .x_share1(d4_P3_23_s1), .y_share0(d4_G3_15_s0), .y_share1(d4_G3_15_s1), .rand(r_t104), .z_share0(d5_t104_s0), .z_share1(d5_t104_s1));
  assign r_t104 = stage5_share0[20];
  and_module u_and_t105_d5 (.clk(clk), .x_share0(d4_P3_24_s0), .x_share1(d4_P3_24_s1), .y_share0(d4_G3_16_s0), .y_share1(d4_G3_16_s1), .rand(r_t105), .z_share0(d5_t105_s0), .z_share1(d5_t105_s1));
  assign r_t105 = stage5_share0[1];
  and_module u_and_t106_d5 (.clk(clk), .x_share0(d4_P3_25_s0), .x_share1(d4_P3_25_s1), .y_share0(d4_G3_17_s0), .y_share1(d4_G3_17_s1), .rand(r_t106), .z_share0(d5_t106_s0), .z_share1(d5_t106_s1));
  assign r_t106 = stage5_share0[5];
  and_module u_and_t107_d5 (.clk(clk), .x_share0(d4_P3_26_s0), .x_share1(d4_P3_26_s1), .y_share0(d4_G3_18_s0), .y_share1(d4_G3_18_s1), .rand(r_t107), .z_share0(d5_t107_s0), .z_share1(d5_t107_s1));
  assign r_t107 = stage5_share0[2];
  and_module u_and_t108_d5 (.clk(clk), .x_share0(d4_P3_27_s0), .x_share1(d4_P3_27_s1), .y_share0(d4_G3_19_s0), .y_share1(d4_G3_19_s1), .rand(r_t108), .z_share0(d5_t108_s0), .z_share1(d5_t108_s1));
  assign r_t108 = stage5_share0[21];
  and_module u_and_t109_d5 (.clk(clk), .x_share0(d4_P3_28_s0), .x_share1(d4_P3_28_s1), .y_share0(d4_G3_20_s0), .y_share1(d4_G3_20_s1), .rand(r_t109), .z_share0(d5_t109_s0), .z_share1(d5_t109_s1));
  assign r_t109 = stage5_share0[0];
  and_module u_and_t110_d5 (.clk(clk), .x_share0(d4_P3_29_s0), .x_share1(d4_P3_29_s1), .y_share0(d4_G3_21_s0), .y_share1(d4_G3_21_s1), .rand(r_t110), .z_share0(d5_t110_s0), .z_share1(d5_t110_s1));
  assign r_t110 = stage5_share0[8];
  and_module u_and_t111_d5 (.clk(clk), .x_share0(d4_P3_30_s0), .x_share1(d4_P3_30_s1), .y_share0(d4_G3_22_s0), .y_share1(d4_G3_22_s1), .rand(r_t111), .z_share0(d5_t111_s0), .z_share1(d5_t111_s1));
  assign r_t111 = stage5_share0[12];
  and_module u_and_t112_d5 (.clk(clk), .x_share0(d4_P3_31_s0), .x_share1(d4_P3_31_s1), .y_share0(d4_G3_23_s0), .y_share1(d4_G3_23_s1), .rand(r_t112), .z_share0(d5_t112_s0), .z_share1(d5_t112_s1));
  assign r_t112 = stage5_share0[2];
  and_module u_and_t113_d5 (.clk(clk), .x_share0(d4_P4_16_s0), .x_share1(d4_P4_16_s1), .y_share0(d4_G0_0_s0), .y_share1(d4_G0_0_s1), .rand(r_t113), .z_share0(d5_t113_s0), .z_share1(d5_t113_s1));
  assign r_t113 = stage5_share0[0];
  and_module u_and_t114_d5 (.clk(clk), .x_share0(d4_P4_17_s0), .x_share1(d4_P4_17_s1), .y_share0(d4_G1_1_s0), .y_share1(d4_G1_1_s1), .rand(r_t114), .z_share0(d5_t114_s0), .z_share1(d5_t114_s1));
  assign r_t114 = stage5_share0[6];
  and_module u_and_t115_d5 (.clk(clk), .x_share0(d4_P4_18_s0), .x_share1(d4_P4_18_s1), .y_share0(d4_G2_2_s0), .y_share1(d4_G2_2_s1), .rand(r_t115), .z_share0(d5_t115_s0), .z_share1(d5_t115_s1));
  assign r_t115 = stage5_share0[7];
  and_module u_and_t116_d5 (.clk(clk), .x_share0(d4_P4_19_s0), .x_share1(d4_P4_19_s1), .y_share0(d4_G2_3_s0), .y_share1(d4_G2_3_s1), .rand(r_t116), .z_share0(d5_t116_s0), .z_share1(d5_t116_s1));
  assign r_t116 = stage5_share0[10];
  and_module u_and_t117_d5 (.clk(clk), .x_share0(d4_P4_20_s0), .x_share1(d4_P4_20_s1), .y_share0(d4_G3_4_s0), .y_share1(d4_G3_4_s1), .rand(r_t117), .z_share0(d5_t117_s0), .z_share1(d5_t117_s1));
  assign r_t117 = stage5_share0[5];
  and_module u_and_t118_d5 (.clk(clk), .x_share0(d4_P4_21_s0), .x_share1(d4_P4_21_s1), .y_share0(d4_G3_5_s0), .y_share1(d4_G3_5_s1), .rand(r_t118), .z_share0(d5_t118_s0), .z_share1(d5_t118_s1));
  assign r_t118 = stage5_share0[12];
  and_module u_and_t119_d5 (.clk(clk), .x_share0(d4_P4_22_s0), .x_share1(d4_P4_22_s1), .y_share0(d4_G3_6_s0), .y_share1(d4_G3_6_s1), .rand(r_t119), .z_share0(d5_t119_s0), .z_share1(d5_t119_s1));
  assign r_t119 = stage5_share0[8];
  and_module u_and_t120_d5 (.clk(clk), .x_share0(d4_P4_23_s0), .x_share1(d4_P4_23_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t120), .z_share0(d5_t120_s0), .z_share1(d5_t120_s1));
  assign r_t120 = stage5_share0[14];
  and_module u_and_t121_d5 (.clk(clk), .x_share0(d4_P4_24_s0), .x_share1(d4_P4_24_s1), .y_share0(d4_G4_8_s0), .y_share1(d4_G4_8_s1), .rand(r_t121), .z_share0(d5_t121_s0), .z_share1(d5_t121_s1));
  assign r_t121 = stage5_share0[21];
  and_module u_and_t122_d5 (.clk(clk), .x_share0(d4_P4_25_s0), .x_share1(d4_P4_25_s1), .y_share0(d4_G4_9_s0), .y_share1(d4_G4_9_s1), .rand(r_t122), .z_share0(d5_t122_s0), .z_share1(d5_t122_s1));
  assign r_t122 = stage5_share0[22];
  and_module u_and_t123_d5 (.clk(clk), .x_share0(d4_P4_26_s0), .x_share1(d4_P4_26_s1), .y_share0(d4_G4_10_s0), .y_share1(d4_G4_10_s1), .rand(r_t123), .z_share0(d5_t123_s0), .z_share1(d5_t123_s1));
  assign r_t123 = stage5_share0[23];
  and_module u_and_t124_d5 (.clk(clk), .x_share0(d4_P4_27_s0), .x_share1(d4_P4_27_s1), .y_share0(d4_G4_11_s0), .y_share1(d4_G4_11_s1), .rand(r_t124), .z_share0(d5_t124_s0), .z_share1(d5_t124_s1));
  assign r_t124 = stage5_share0[18];
  and_module u_and_t125_d5 (.clk(clk), .x_share0(d4_P4_28_s0), .x_share1(d4_P4_28_s1), .y_share0(d4_G4_12_s0), .y_share1(d4_G4_12_s1), .rand(r_t125), .z_share0(d5_t125_s0), .z_share1(d5_t125_s1));
  assign r_t125 = stage5_share0[25];
  and_module u_and_t126_d5 (.clk(clk), .x_share0(d4_P4_29_s0), .x_share1(d4_P4_29_s1), .y_share0(d4_G4_13_s0), .y_share1(d4_G4_13_s1), .rand(r_t126), .z_share0(d5_t126_s0), .z_share1(d5_t126_s1));
  assign r_t126 = stage5_share0[26];
  and_module u_and_t127_d5 (.clk(clk), .x_share0(d4_P4_30_s0), .x_share1(d4_P4_30_s1), .y_share0(d4_G4_14_s0), .y_share1(d4_G4_14_s1), .rand(r_t127), .z_share0(d5_t127_s0), .z_share1(d5_t127_s1));
  assign r_t127 = stage5_share0[25];
  and_module u_and_t96_d5 (.clk(clk), .x_share0(d4_P3_15_s0), .x_share1(d4_P3_15_s1), .y_share0(d4_G3_7_s0), .y_share1(d4_G3_7_s1), .rand(r_t96), .z_share0(d5_t96_s0), .z_share1(d5_t96_s1));
  assign r_t96 = stage5_share0[6];
  and_module u_and_t97_d5 (.clk(clk), .x_share0(d4_P3_16_s0), .x_share1(d4_P3_16_s1), .y_share0(d4_G3_8_s0), .y_share1(d4_G3_8_s1), .rand(r_t97), .z_share0(d5_t97_s0), .z_share1(d5_t97_s1));
  assign r_t97 = stage5_share0[2];
  and_module u_and_t98_d5 (.clk(clk), .x_share0(d4_P3_17_s0), .x_share1(d4_P3_17_s1), .y_share0(d4_G3_9_s0), .y_share1(d4_G3_9_s1), .rand(r_t98), .z_share0(d5_t98_s0), .z_share1(d5_t98_s1));
  assign r_t98 = stage5_share0[7];
  and_module u_and_t99_d5 (.clk(clk), .x_share0(d4_P3_18_s0), .x_share1(d4_P3_18_s1), .y_share0(d4_G3_10_s0), .y_share1(d4_G3_10_s1), .rand(r_t99), .z_share0(d5_t99_s0), .z_share1(d5_t99_s1));
  assign r_t99 = stage5_share0[12];
  reg_module u_reg_G4_31_d6 (.clk(clk), .input_share0(d5_G4_31_s0), .input_share1(d5_G4_31_s1), .output_share0(d6_G4_31_s0), .output_share1(d6_G4_31_s1));
  xor_module u_xor_G5_31_d6 (.x_share0(d6_t128_s0), .x_share1(d6_t128_s1), .y_share0(d6_G4_31_s0), .y_share1(d6_G4_31_s1), .z_share0(d6_G5_31_s0), .z_share1(d6_G5_31_s1));
  and_module u_and_t128_d6 (.clk(clk), .x_share0(d5_P4_31_s0), .x_share1(d5_P4_31_s1), .y_share0(d5_G4_15_s0), .y_share1(d5_G4_15_s1), .rand(r_t128), .z_share0(d6_t128_s0), .z_share1(d6_t128_s1));
  assign r_t128 = stage6_share0[9];

  // Output assignments
  assign o_share0[0] = d0_o0_s0;
  assign o_share1[0] = d0_o0_s1;
  assign o_share0[1] = d1_o1_s0;
  assign o_share1[1] = d1_o1_s1;
  assign o_share0[2] = d2_o2_s0;
  assign o_share1[2] = d2_o2_s1;
  assign o_share0[3] = d2_o3_s0;
  assign o_share1[3] = d2_o3_s1;
  assign o_share0[4] = d3_o4_s0;
  assign o_share1[4] = d3_o4_s1;
  assign o_share0[5] = d3_o5_s0;
  assign o_share1[5] = d3_o5_s1;
  assign o_share0[6] = d3_o6_s0;
  assign o_share1[6] = d3_o6_s1;
  assign o_share0[7] = d3_o7_s0;
  assign o_share1[7] = d3_o7_s1;
  assign o_share0[8] = d4_o8_s0;
  assign o_share1[8] = d4_o8_s1;
  assign o_share0[9] = d4_o9_s0;
  assign o_share1[9] = d4_o9_s1;
  assign o_share0[10] = d4_o10_s0;
  assign o_share1[10] = d4_o10_s1;
  assign o_share0[11] = d4_o11_s0;
  assign o_share1[11] = d4_o11_s1;
  assign o_share0[12] = d4_o12_s0;
  assign o_share1[12] = d4_o12_s1;
  assign o_share0[13] = d4_o13_s0;
  assign o_share1[13] = d4_o13_s1;
  assign o_share0[14] = d4_o14_s0;
  assign o_share1[14] = d4_o14_s1;
  assign o_share0[15] = d4_o15_s0;
  assign o_share1[15] = d4_o15_s1;
  assign o_share0[16] = d5_o16_s0;
  assign o_share1[16] = d5_o16_s1;
  assign o_share0[17] = d5_o17_s0;
  assign o_share1[17] = d5_o17_s1;
  assign o_share0[18] = d5_o18_s0;
  assign o_share1[18] = d5_o18_s1;
  assign o_share0[19] = d5_o19_s0;
  assign o_share1[19] = d5_o19_s1;
  assign o_share0[20] = d5_o20_s0;
  assign o_share1[20] = d5_o20_s1;
  assign o_share0[21] = d5_o21_s0;
  assign o_share1[21] = d5_o21_s1;
  assign o_share0[22] = d5_o22_s0;
  assign o_share1[22] = d5_o22_s1;
  assign o_share0[23] = d5_o23_s0;
  assign o_share1[23] = d5_o23_s1;
  assign o_share0[24] = d5_o24_s0;
  assign o_share1[24] = d5_o24_s1;
  assign o_share0[25] = d5_o25_s0;
  assign o_share1[25] = d5_o25_s1;
  assign o_share0[26] = d5_o26_s0;
  assign o_share1[26] = d5_o26_s1;
  assign o_share0[27] = d5_o27_s0;
  assign o_share1[27] = d5_o27_s1;
  assign o_share0[28] = d5_o28_s0;
  assign o_share1[28] = d5_o28_s1;
  assign o_share0[29] = d5_o29_s0;
  assign o_share1[29] = d5_o29_s1;
  assign o_share0[30] = d5_o30_s0;
  assign o_share1[30] = d5_o30_s1;
  assign o_share0[31] = d5_o31_s0;
  assign o_share1[31] = d5_o31_s1;

endmodule
